package flowtest;
import FIFO::*;
import FIFOF::*;
import datatypes::*;
import SpecialFIFOs:: * ;
import Real::*;
import Vector::*;
import compact::*;


#define L0 128 
(*synthesize*)
module mkFlowTest();

CompactTree px <- mkCompactTree;
	rule push_data;
	Vector#(L0,Int#(16)) r = newVector;
		r[0]=27;
		r[1]=0;
		r[2]=96;
		r[3]=0;
		r[4]=32;
		r[5]=95;
		r[6]=34;
		r[7]=0;
		r[8]=190;
		r[9]=0;
		r[10]=0;
		r[11]=0;
		r[12]=0;
		r[13]=0;
		r[14]=0;
		r[15]=0;
		r[16]=0;
		r[17]=0;
		r[18]=0;
		r[19]=0;
		r[20]=20;
		r[21]=0;
		r[22]=0;
		r[23]=180;
		r[24]=0;
		r[25]=13;
		r[26]=25;
		r[27]=194;
		r[28]=0;
		r[29]=0;
		r[30]=195;
		r[31]=105;
		r[32]=0;
		r[33]=182;
		r[34]=55;
		r[35]=16;
		r[36]=0;
		r[37]=0;
		r[38]=0;
		r[39]=42;
		r[40]=0;
		r[41]=0;
		r[42]=0;
		r[43]=72;
		r[44]=64;
		r[45]=101;
		r[46]=0;
		r[47]=80;
		r[48]=137;
		r[49]=140;
		r[50]=56;
		r[51]=24;
		r[52]=0;
		r[53]=114;
		r[54]=0;
		r[55]=0;
		r[56]=0;
		r[57]=0;
		r[58]=110;
		r[59]=187;
		r[60]=169;
		r[61]=137;
		r[62]=47;
		r[63]=163;
		r[64]=62;
		r[65]=161;
		r[66]=72;
		r[67]=0;
		r[68]=0;
		r[69]=161;
		r[70]=132;
		r[71]=0;
		r[72]=66;
		r[73]=0;
		r[74]=86;
		r[75]=106;
		r[76]=48;
		r[77]=178;
		r[78]=19;
		r[79]=0;
		r[80]=0;
		r[81]=88;
		r[82]=0;
		r[83]=0;
		r[84]=0;
		r[85]=0;
		r[86]=0;
		r[87]=0;
		r[88]=0;
		r[89]=0;
		r[90]=13;
		r[91]=40;
		r[92]=0;
		r[93]=54;
		r[94]=70;
		r[95]=151;
		r[96]=65;
		r[97]=0;
		r[98]=40;
		r[99]=30;
		r[100]=0;
		r[101]=0;
		r[102]=151;
		r[103]=58;
		r[104]=0;
		r[105]=19;
		r[106]=64;
		r[107]=68;
		r[108]=0;
		r[109]=126;
		r[110]=126;
		r[111]=0;
		r[112]=0;
		r[113]=147;
		r[114]=122;
		r[115]=0;
		r[116]=0;
		r[117]=23;
		r[118]=0;
		r[119]=199;
		r[120]=0;
		r[121]=100;
		r[122]=0;
		r[123]=0;
		r[124]=132;
		r[125]=134;
		r[126]=0;
		r[127]=168;
	px.put(unpack(pack(r)));
	endrule
	rule get_data;
	let d <- px.get;
	Vector#(L0, Int#(16)) dx = unpack(d);
	for(int i=0; i<L0; i=i+1)
	$display("%d",dx[i]);
	$finish(0);
	endrule
endmodule
endpackage