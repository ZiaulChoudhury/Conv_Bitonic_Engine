package bitonic;
import FIFO::*;
import FIFOF::*;
import datatypes::*;
import SpecialFIFOs:: * ;
import Real::*;
import Vector::*;
#define L0 256

interface Bitonic;
        method Action put(Vector#(L0, Int#(32)) datas);
        method ActionValue#(Vector#(L0, Int#(32))) get;
endinterface


function Vector#(2,Int#(32)) min_max(Bit#(32) pkt1, Bit#(32) pkt2);
	Int#(8)  p1_partition = unpack(pkt1[7:0]);
	Int#(8)  p2_partition = unpack(pkt2[7:0]);
	Int#(8)  p1_conv      = unpack(pkt1[15:8]);
	Int#(8)  p2_conv      = unpack(pkt2[15:8]);
	Vector#(2,Int#(32)) sort = newVector;
	if (p1_partition < p2_partition || (p1_partition == p2_partition && p1_conv < p2_conv)) begin
		 sort[0] = unpack(pkt1); sort[1] = unpack(pkt2); end
	else begin
		 sort[1] = unpack(pkt1); sort[0] = unpack(pkt2); end
	return sort;
endfunction


(*synthesize*)
module mkBitonic(Bitonic);
Reg#(Int#(32)) s0[L0];
Reg#(Int#(32)) s1[L0];
Reg#(Int#(32)) s2[L0];
Reg#(Int#(32)) s3[L0];
Reg#(Int#(32)) s4[L0];
Reg#(Int#(32)) s5[L0];
Reg#(Int#(32)) s6[L0];
Reg#(Int#(32)) s7[L0];
Reg#(Int#(32)) s8[L0];
Reg#(Int#(32)) s9[L0];
Reg#(Int#(32)) s10[L0];
Reg#(Int#(32)) s11[L0];
Reg#(Int#(32)) s12[L0];
Reg#(Int#(32)) s13[L0];
Reg#(Int#(32)) s14[L0];
Reg#(Int#(32)) s15[L0];
Reg#(Int#(32)) s16[L0];
Reg#(Int#(32)) s17[L0];
Reg#(Int#(32)) s18[L0];
Reg#(Int#(32)) s19[L0];
Reg#(Int#(32)) s20[L0];
Reg#(Int#(32)) s21[L0];
Reg#(Int#(32)) s22[L0];
Reg#(Int#(32)) s23[L0];
Reg#(Int#(32)) s24[L0];
Reg#(Int#(32)) s25[L0];
Reg#(Int#(32)) s26[L0];
Reg#(Int#(32)) s27[L0];
Reg#(Int#(32)) s28[L0];
Reg#(Int#(32)) s29[L0];
Reg#(Int#(32)) s30[L0];
Reg#(Int#(32)) s31[L0];
Reg#(Int#(32)) s32[L0];
Reg#(Int#(32)) s33[L0];
Reg#(Int#(32)) s34[L0];
Reg#(Int#(32)) s35[L0];
Reg#(Int#(32)) s36[L0];

for(int i =0; i<L0; i = i + 1) begin
s0[i] <- mkReg(0);
s1[i] <- mkReg(0);
s2[i] <- mkReg(0);
s3[i] <- mkReg(0);
s4[i] <- mkReg(0);
s5[i] <- mkReg(0);
s6[i] <- mkReg(0);
s7[i] <- mkReg(0);
s8[i] <- mkReg(0);
s9[i] <- mkReg(0);
s10[i] <- mkReg(0);
s11[i] <- mkReg(0);
s12[i] <- mkReg(0);
s13[i] <- mkReg(0);
s14[i] <- mkReg(0);
s15[i] <- mkReg(0);
s16[i] <- mkReg(0);
s17[i] <- mkReg(0);
s18[i] <- mkReg(0);
s19[i] <- mkReg(0);
s20[i] <- mkReg(0);
s21[i] <- mkReg(0);
s22[i] <- mkReg(0);
s23[i] <- mkReg(0);
s24[i] <- mkReg(0);
s25[i] <- mkReg(0);
s26[i] <- mkReg(0);
s27[i] <- mkReg(0);
s28[i] <- mkReg(0);
s29[i] <- mkReg(0);
s30[i] <- mkReg(0);
s31[i] <- mkReg(0);
s32[i] <- mkReg(0);
s33[i] <- mkReg(0);
s34[i] <- mkReg(0);
s35[i] <- mkReg(0);
s36[i] <- mkReg(0);
end
FIFOF#(Bit#(1)) p0 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p1 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p2 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p3 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p4 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p5 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p6 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p7 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p8 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p9 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p10 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p11 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p12 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p13 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p14 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p15 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p16 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p17 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p18 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p19 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p20 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p21 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p22 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p23 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p24 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p25 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p26 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p27 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p28 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p29 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p30 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p31 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p32 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p33 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p34 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p35 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p36 <- mkPipelineFIFOF;
rule _Q01;
	p0.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S1i0 = min_max(pack(s0[mod*i+0]) , pack(s0[mod*i+0+mod/2]));
		if ((i/1)%2 == 0) begin
			s1[mod*i+0] <= _S1i0[0];
			s1[mod*i+0+mod/2] <= _S1i0[1];
		end
		else begin
			s1[mod*i+0] <= _S1i0[1];
			s1[mod*i+0+mod/2] <= _S1i0[0];
		end
	end
	p1.enq(1);
endrule
rule _Q12;
	p1.deq;
	let mod = 4;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S2i0 = min_max(pack(s1[mod*i+0]) , pack(s1[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S2i1 = min_max(pack(s1[mod*i+1]) , pack(s1[mod*i+1+mod/2]));
		if ((i/1)%2 == 0) begin
			s2[mod*i+0] <= _S2i0[0];
			s2[mod*i+0+mod/2] <= _S2i0[1];
			s2[mod*i+1] <= _S2i1[0];
			s2[mod*i+1+mod/2] <= _S2i1[1];
		end
		else begin
			s2[mod*i+0] <= _S2i0[1];
			s2[mod*i+0+mod/2] <= _S2i0[0];
			s2[mod*i+1] <= _S2i1[1];
			s2[mod*i+1+mod/2] <= _S2i1[0];
		end
	end
	p2.enq(1);
endrule
rule _Q11;
	p2.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S3i0 = min_max(pack(s2[mod*i+0]) , pack(s2[mod*i+0+mod/2]));
		if ((i/2)%2 == 0) begin
			s3[mod*i+0] <= _S3i0[0];
			s3[mod*i+0+mod/2] <= _S3i0[1];
		end
		else begin
			s3[mod*i+0] <= _S3i0[1];
			s3[mod*i+0+mod/2] <= _S3i0[0];
		end
	end
	p3.enq(1);
endrule
rule _Q23;
	p3.deq;
	let mod = 8;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S4i0 = min_max(pack(s3[mod*i+0]) , pack(s3[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S4i1 = min_max(pack(s3[mod*i+1]) , pack(s3[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S4i2 = min_max(pack(s3[mod*i+2]) , pack(s3[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S4i3 = min_max(pack(s3[mod*i+3]) , pack(s3[mod*i+3+mod/2]));
		if ((i/1)%2 == 0) begin
			s4[mod*i+0] <= _S4i0[0];
			s4[mod*i+0+mod/2] <= _S4i0[1];
			s4[mod*i+1] <= _S4i1[0];
			s4[mod*i+1+mod/2] <= _S4i1[1];
			s4[mod*i+2] <= _S4i2[0];
			s4[mod*i+2+mod/2] <= _S4i2[1];
			s4[mod*i+3] <= _S4i3[0];
			s4[mod*i+3+mod/2] <= _S4i3[1];
		end
		else begin
			s4[mod*i+0] <= _S4i0[1];
			s4[mod*i+0+mod/2] <= _S4i0[0];
			s4[mod*i+1] <= _S4i1[1];
			s4[mod*i+1+mod/2] <= _S4i1[0];
			s4[mod*i+2] <= _S4i2[1];
			s4[mod*i+2+mod/2] <= _S4i2[0];
			s4[mod*i+3] <= _S4i3[1];
			s4[mod*i+3+mod/2] <= _S4i3[0];
		end
	end
	p4.enq(1);
endrule
rule _Q22;
	p4.deq;
	let mod = 4;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S5i0 = min_max(pack(s4[mod*i+0]) , pack(s4[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S5i1 = min_max(pack(s4[mod*i+1]) , pack(s4[mod*i+1+mod/2]));
		if ((i/2)%2 == 0) begin
			s5[mod*i+0] <= _S5i0[0];
			s5[mod*i+0+mod/2] <= _S5i0[1];
			s5[mod*i+1] <= _S5i1[0];
			s5[mod*i+1+mod/2] <= _S5i1[1];
		end
		else begin
			s5[mod*i+0] <= _S5i0[1];
			s5[mod*i+0+mod/2] <= _S5i0[0];
			s5[mod*i+1] <= _S5i1[1];
			s5[mod*i+1+mod/2] <= _S5i1[0];
		end
	end
	p5.enq(1);
endrule
rule _Q21;
	p5.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S6i0 = min_max(pack(s5[mod*i+0]) , pack(s5[mod*i+0+mod/2]));
		if ((i/4)%2 == 0) begin
			s6[mod*i+0] <= _S6i0[0];
			s6[mod*i+0+mod/2] <= _S6i0[1];
		end
		else begin
			s6[mod*i+0] <= _S6i0[1];
			s6[mod*i+0+mod/2] <= _S6i0[0];
		end
	end
	p6.enq(1);
endrule
rule _Q34;
	p6.deq;
	let mod = 16;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S7i0 = min_max(pack(s6[mod*i+0]) , pack(s6[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S7i1 = min_max(pack(s6[mod*i+1]) , pack(s6[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S7i2 = min_max(pack(s6[mod*i+2]) , pack(s6[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S7i3 = min_max(pack(s6[mod*i+3]) , pack(s6[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S7i4 = min_max(pack(s6[mod*i+4]) , pack(s6[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S7i5 = min_max(pack(s6[mod*i+5]) , pack(s6[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S7i6 = min_max(pack(s6[mod*i+6]) , pack(s6[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S7i7 = min_max(pack(s6[mod*i+7]) , pack(s6[mod*i+7+mod/2]));
		if ((i/1)%2 == 0) begin
			s7[mod*i+0] <= _S7i0[0];
			s7[mod*i+0+mod/2] <= _S7i0[1];
			s7[mod*i+1] <= _S7i1[0];
			s7[mod*i+1+mod/2] <= _S7i1[1];
			s7[mod*i+2] <= _S7i2[0];
			s7[mod*i+2+mod/2] <= _S7i2[1];
			s7[mod*i+3] <= _S7i3[0];
			s7[mod*i+3+mod/2] <= _S7i3[1];
			s7[mod*i+4] <= _S7i4[0];
			s7[mod*i+4+mod/2] <= _S7i4[1];
			s7[mod*i+5] <= _S7i5[0];
			s7[mod*i+5+mod/2] <= _S7i5[1];
			s7[mod*i+6] <= _S7i6[0];
			s7[mod*i+6+mod/2] <= _S7i6[1];
			s7[mod*i+7] <= _S7i7[0];
			s7[mod*i+7+mod/2] <= _S7i7[1];
		end
		else begin
			s7[mod*i+0] <= _S7i0[1];
			s7[mod*i+0+mod/2] <= _S7i0[0];
			s7[mod*i+1] <= _S7i1[1];
			s7[mod*i+1+mod/2] <= _S7i1[0];
			s7[mod*i+2] <= _S7i2[1];
			s7[mod*i+2+mod/2] <= _S7i2[0];
			s7[mod*i+3] <= _S7i3[1];
			s7[mod*i+3+mod/2] <= _S7i3[0];
			s7[mod*i+4] <= _S7i4[1];
			s7[mod*i+4+mod/2] <= _S7i4[0];
			s7[mod*i+5] <= _S7i5[1];
			s7[mod*i+5+mod/2] <= _S7i5[0];
			s7[mod*i+6] <= _S7i6[1];
			s7[mod*i+6+mod/2] <= _S7i6[0];
			s7[mod*i+7] <= _S7i7[1];
			s7[mod*i+7+mod/2] <= _S7i7[0];
		end
	end
	p7.enq(1);
endrule
rule _Q33;
	p7.deq;
	let mod = 8;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S8i0 = min_max(pack(s7[mod*i+0]) , pack(s7[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S8i1 = min_max(pack(s7[mod*i+1]) , pack(s7[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S8i2 = min_max(pack(s7[mod*i+2]) , pack(s7[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S8i3 = min_max(pack(s7[mod*i+3]) , pack(s7[mod*i+3+mod/2]));
		if ((i/2)%2 == 0) begin
			s8[mod*i+0] <= _S8i0[0];
			s8[mod*i+0+mod/2] <= _S8i0[1];
			s8[mod*i+1] <= _S8i1[0];
			s8[mod*i+1+mod/2] <= _S8i1[1];
			s8[mod*i+2] <= _S8i2[0];
			s8[mod*i+2+mod/2] <= _S8i2[1];
			s8[mod*i+3] <= _S8i3[0];
			s8[mod*i+3+mod/2] <= _S8i3[1];
		end
		else begin
			s8[mod*i+0] <= _S8i0[1];
			s8[mod*i+0+mod/2] <= _S8i0[0];
			s8[mod*i+1] <= _S8i1[1];
			s8[mod*i+1+mod/2] <= _S8i1[0];
			s8[mod*i+2] <= _S8i2[1];
			s8[mod*i+2+mod/2] <= _S8i2[0];
			s8[mod*i+3] <= _S8i3[1];
			s8[mod*i+3+mod/2] <= _S8i3[0];
		end
	end
	p8.enq(1);
endrule
rule _Q32;
	p8.deq;
	let mod = 4;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S9i0 = min_max(pack(s8[mod*i+0]) , pack(s8[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S9i1 = min_max(pack(s8[mod*i+1]) , pack(s8[mod*i+1+mod/2]));
		if ((i/4)%2 == 0) begin
			s9[mod*i+0] <= _S9i0[0];
			s9[mod*i+0+mod/2] <= _S9i0[1];
			s9[mod*i+1] <= _S9i1[0];
			s9[mod*i+1+mod/2] <= _S9i1[1];
		end
		else begin
			s9[mod*i+0] <= _S9i0[1];
			s9[mod*i+0+mod/2] <= _S9i0[0];
			s9[mod*i+1] <= _S9i1[1];
			s9[mod*i+1+mod/2] <= _S9i1[0];
		end
	end
	p9.enq(1);
endrule
rule _Q31;
	p9.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S10i0 = min_max(pack(s9[mod*i+0]) , pack(s9[mod*i+0+mod/2]));
		if ((i/8)%2 == 0) begin
			s10[mod*i+0] <= _S10i0[0];
			s10[mod*i+0+mod/2] <= _S10i0[1];
		end
		else begin
			s10[mod*i+0] <= _S10i0[1];
			s10[mod*i+0+mod/2] <= _S10i0[0];
		end
	end
	p10.enq(1);
endrule
rule _Q45;
	p10.deq;
	let mod = 32;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S11i0 = min_max(pack(s10[mod*i+0]) , pack(s10[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S11i1 = min_max(pack(s10[mod*i+1]) , pack(s10[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S11i2 = min_max(pack(s10[mod*i+2]) , pack(s10[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S11i3 = min_max(pack(s10[mod*i+3]) , pack(s10[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S11i4 = min_max(pack(s10[mod*i+4]) , pack(s10[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S11i5 = min_max(pack(s10[mod*i+5]) , pack(s10[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S11i6 = min_max(pack(s10[mod*i+6]) , pack(s10[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S11i7 = min_max(pack(s10[mod*i+7]) , pack(s10[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S11i8 = min_max(pack(s10[mod*i+8]) , pack(s10[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S11i9 = min_max(pack(s10[mod*i+9]) , pack(s10[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S11i10 = min_max(pack(s10[mod*i+10]) , pack(s10[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S11i11 = min_max(pack(s10[mod*i+11]) , pack(s10[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S11i12 = min_max(pack(s10[mod*i+12]) , pack(s10[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S11i13 = min_max(pack(s10[mod*i+13]) , pack(s10[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S11i14 = min_max(pack(s10[mod*i+14]) , pack(s10[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S11i15 = min_max(pack(s10[mod*i+15]) , pack(s10[mod*i+15+mod/2]));
		if ((i/1)%2 == 0) begin
			s11[mod*i+0] <= _S11i0[0];
			s11[mod*i+0+mod/2] <= _S11i0[1];
			s11[mod*i+1] <= _S11i1[0];
			s11[mod*i+1+mod/2] <= _S11i1[1];
			s11[mod*i+2] <= _S11i2[0];
			s11[mod*i+2+mod/2] <= _S11i2[1];
			s11[mod*i+3] <= _S11i3[0];
			s11[mod*i+3+mod/2] <= _S11i3[1];
			s11[mod*i+4] <= _S11i4[0];
			s11[mod*i+4+mod/2] <= _S11i4[1];
			s11[mod*i+5] <= _S11i5[0];
			s11[mod*i+5+mod/2] <= _S11i5[1];
			s11[mod*i+6] <= _S11i6[0];
			s11[mod*i+6+mod/2] <= _S11i6[1];
			s11[mod*i+7] <= _S11i7[0];
			s11[mod*i+7+mod/2] <= _S11i7[1];
			s11[mod*i+8] <= _S11i8[0];
			s11[mod*i+8+mod/2] <= _S11i8[1];
			s11[mod*i+9] <= _S11i9[0];
			s11[mod*i+9+mod/2] <= _S11i9[1];
			s11[mod*i+10] <= _S11i10[0];
			s11[mod*i+10+mod/2] <= _S11i10[1];
			s11[mod*i+11] <= _S11i11[0];
			s11[mod*i+11+mod/2] <= _S11i11[1];
			s11[mod*i+12] <= _S11i12[0];
			s11[mod*i+12+mod/2] <= _S11i12[1];
			s11[mod*i+13] <= _S11i13[0];
			s11[mod*i+13+mod/2] <= _S11i13[1];
			s11[mod*i+14] <= _S11i14[0];
			s11[mod*i+14+mod/2] <= _S11i14[1];
			s11[mod*i+15] <= _S11i15[0];
			s11[mod*i+15+mod/2] <= _S11i15[1];
		end
		else begin
			s11[mod*i+0] <= _S11i0[1];
			s11[mod*i+0+mod/2] <= _S11i0[0];
			s11[mod*i+1] <= _S11i1[1];
			s11[mod*i+1+mod/2] <= _S11i1[0];
			s11[mod*i+2] <= _S11i2[1];
			s11[mod*i+2+mod/2] <= _S11i2[0];
			s11[mod*i+3] <= _S11i3[1];
			s11[mod*i+3+mod/2] <= _S11i3[0];
			s11[mod*i+4] <= _S11i4[1];
			s11[mod*i+4+mod/2] <= _S11i4[0];
			s11[mod*i+5] <= _S11i5[1];
			s11[mod*i+5+mod/2] <= _S11i5[0];
			s11[mod*i+6] <= _S11i6[1];
			s11[mod*i+6+mod/2] <= _S11i6[0];
			s11[mod*i+7] <= _S11i7[1];
			s11[mod*i+7+mod/2] <= _S11i7[0];
			s11[mod*i+8] <= _S11i8[1];
			s11[mod*i+8+mod/2] <= _S11i8[0];
			s11[mod*i+9] <= _S11i9[1];
			s11[mod*i+9+mod/2] <= _S11i9[0];
			s11[mod*i+10] <= _S11i10[1];
			s11[mod*i+10+mod/2] <= _S11i10[0];
			s11[mod*i+11] <= _S11i11[1];
			s11[mod*i+11+mod/2] <= _S11i11[0];
			s11[mod*i+12] <= _S11i12[1];
			s11[mod*i+12+mod/2] <= _S11i12[0];
			s11[mod*i+13] <= _S11i13[1];
			s11[mod*i+13+mod/2] <= _S11i13[0];
			s11[mod*i+14] <= _S11i14[1];
			s11[mod*i+14+mod/2] <= _S11i14[0];
			s11[mod*i+15] <= _S11i15[1];
			s11[mod*i+15+mod/2] <= _S11i15[0];
		end
	end
	p11.enq(1);
endrule
rule _Q44;
	p11.deq;
	let mod = 16;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S12i0 = min_max(pack(s11[mod*i+0]) , pack(s11[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S12i1 = min_max(pack(s11[mod*i+1]) , pack(s11[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S12i2 = min_max(pack(s11[mod*i+2]) , pack(s11[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S12i3 = min_max(pack(s11[mod*i+3]) , pack(s11[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S12i4 = min_max(pack(s11[mod*i+4]) , pack(s11[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S12i5 = min_max(pack(s11[mod*i+5]) , pack(s11[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S12i6 = min_max(pack(s11[mod*i+6]) , pack(s11[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S12i7 = min_max(pack(s11[mod*i+7]) , pack(s11[mod*i+7+mod/2]));
		if ((i/2)%2 == 0) begin
			s12[mod*i+0] <= _S12i0[0];
			s12[mod*i+0+mod/2] <= _S12i0[1];
			s12[mod*i+1] <= _S12i1[0];
			s12[mod*i+1+mod/2] <= _S12i1[1];
			s12[mod*i+2] <= _S12i2[0];
			s12[mod*i+2+mod/2] <= _S12i2[1];
			s12[mod*i+3] <= _S12i3[0];
			s12[mod*i+3+mod/2] <= _S12i3[1];
			s12[mod*i+4] <= _S12i4[0];
			s12[mod*i+4+mod/2] <= _S12i4[1];
			s12[mod*i+5] <= _S12i5[0];
			s12[mod*i+5+mod/2] <= _S12i5[1];
			s12[mod*i+6] <= _S12i6[0];
			s12[mod*i+6+mod/2] <= _S12i6[1];
			s12[mod*i+7] <= _S12i7[0];
			s12[mod*i+7+mod/2] <= _S12i7[1];
		end
		else begin
			s12[mod*i+0] <= _S12i0[1];
			s12[mod*i+0+mod/2] <= _S12i0[0];
			s12[mod*i+1] <= _S12i1[1];
			s12[mod*i+1+mod/2] <= _S12i1[0];
			s12[mod*i+2] <= _S12i2[1];
			s12[mod*i+2+mod/2] <= _S12i2[0];
			s12[mod*i+3] <= _S12i3[1];
			s12[mod*i+3+mod/2] <= _S12i3[0];
			s12[mod*i+4] <= _S12i4[1];
			s12[mod*i+4+mod/2] <= _S12i4[0];
			s12[mod*i+5] <= _S12i5[1];
			s12[mod*i+5+mod/2] <= _S12i5[0];
			s12[mod*i+6] <= _S12i6[1];
			s12[mod*i+6+mod/2] <= _S12i6[0];
			s12[mod*i+7] <= _S12i7[1];
			s12[mod*i+7+mod/2] <= _S12i7[0];
		end
	end
	p12.enq(1);
endrule
rule _Q43;
	p12.deq;
	let mod = 8;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S13i0 = min_max(pack(s12[mod*i+0]) , pack(s12[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S13i1 = min_max(pack(s12[mod*i+1]) , pack(s12[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S13i2 = min_max(pack(s12[mod*i+2]) , pack(s12[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S13i3 = min_max(pack(s12[mod*i+3]) , pack(s12[mod*i+3+mod/2]));
		if ((i/4)%2 == 0) begin
			s13[mod*i+0] <= _S13i0[0];
			s13[mod*i+0+mod/2] <= _S13i0[1];
			s13[mod*i+1] <= _S13i1[0];
			s13[mod*i+1+mod/2] <= _S13i1[1];
			s13[mod*i+2] <= _S13i2[0];
			s13[mod*i+2+mod/2] <= _S13i2[1];
			s13[mod*i+3] <= _S13i3[0];
			s13[mod*i+3+mod/2] <= _S13i3[1];
		end
		else begin
			s13[mod*i+0] <= _S13i0[1];
			s13[mod*i+0+mod/2] <= _S13i0[0];
			s13[mod*i+1] <= _S13i1[1];
			s13[mod*i+1+mod/2] <= _S13i1[0];
			s13[mod*i+2] <= _S13i2[1];
			s13[mod*i+2+mod/2] <= _S13i2[0];
			s13[mod*i+3] <= _S13i3[1];
			s13[mod*i+3+mod/2] <= _S13i3[0];
		end
	end
	p13.enq(1);
endrule
rule _Q42;
	p13.deq;
	let mod = 4;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S14i0 = min_max(pack(s13[mod*i+0]) , pack(s13[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S14i1 = min_max(pack(s13[mod*i+1]) , pack(s13[mod*i+1+mod/2]));
		if ((i/8)%2 == 0) begin
			s14[mod*i+0] <= _S14i0[0];
			s14[mod*i+0+mod/2] <= _S14i0[1];
			s14[mod*i+1] <= _S14i1[0];
			s14[mod*i+1+mod/2] <= _S14i1[1];
		end
		else begin
			s14[mod*i+0] <= _S14i0[1];
			s14[mod*i+0+mod/2] <= _S14i0[0];
			s14[mod*i+1] <= _S14i1[1];
			s14[mod*i+1+mod/2] <= _S14i1[0];
		end
	end
	p14.enq(1);
endrule
rule _Q41;
	p14.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S15i0 = min_max(pack(s14[mod*i+0]) , pack(s14[mod*i+0+mod/2]));
		if ((i/16)%2 == 0) begin
			s15[mod*i+0] <= _S15i0[0];
			s15[mod*i+0+mod/2] <= _S15i0[1];
		end
		else begin
			s15[mod*i+0] <= _S15i0[1];
			s15[mod*i+0+mod/2] <= _S15i0[0];
		end
	end
	p15.enq(1);
endrule
rule _Q56;
	p15.deq;
	let mod = 64;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S16i0 = min_max(pack(s15[mod*i+0]) , pack(s15[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S16i1 = min_max(pack(s15[mod*i+1]) , pack(s15[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S16i2 = min_max(pack(s15[mod*i+2]) , pack(s15[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S16i3 = min_max(pack(s15[mod*i+3]) , pack(s15[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S16i4 = min_max(pack(s15[mod*i+4]) , pack(s15[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S16i5 = min_max(pack(s15[mod*i+5]) , pack(s15[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S16i6 = min_max(pack(s15[mod*i+6]) , pack(s15[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S16i7 = min_max(pack(s15[mod*i+7]) , pack(s15[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S16i8 = min_max(pack(s15[mod*i+8]) , pack(s15[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S16i9 = min_max(pack(s15[mod*i+9]) , pack(s15[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S16i10 = min_max(pack(s15[mod*i+10]) , pack(s15[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S16i11 = min_max(pack(s15[mod*i+11]) , pack(s15[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S16i12 = min_max(pack(s15[mod*i+12]) , pack(s15[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S16i13 = min_max(pack(s15[mod*i+13]) , pack(s15[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S16i14 = min_max(pack(s15[mod*i+14]) , pack(s15[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S16i15 = min_max(pack(s15[mod*i+15]) , pack(s15[mod*i+15+mod/2]));
			 Vector#(2, Int#(32)) _S16i16 = min_max(pack(s15[mod*i+16]) , pack(s15[mod*i+16+mod/2]));
			 Vector#(2, Int#(32)) _S16i17 = min_max(pack(s15[mod*i+17]) , pack(s15[mod*i+17+mod/2]));
			 Vector#(2, Int#(32)) _S16i18 = min_max(pack(s15[mod*i+18]) , pack(s15[mod*i+18+mod/2]));
			 Vector#(2, Int#(32)) _S16i19 = min_max(pack(s15[mod*i+19]) , pack(s15[mod*i+19+mod/2]));
			 Vector#(2, Int#(32)) _S16i20 = min_max(pack(s15[mod*i+20]) , pack(s15[mod*i+20+mod/2]));
			 Vector#(2, Int#(32)) _S16i21 = min_max(pack(s15[mod*i+21]) , pack(s15[mod*i+21+mod/2]));
			 Vector#(2, Int#(32)) _S16i22 = min_max(pack(s15[mod*i+22]) , pack(s15[mod*i+22+mod/2]));
			 Vector#(2, Int#(32)) _S16i23 = min_max(pack(s15[mod*i+23]) , pack(s15[mod*i+23+mod/2]));
			 Vector#(2, Int#(32)) _S16i24 = min_max(pack(s15[mod*i+24]) , pack(s15[mod*i+24+mod/2]));
			 Vector#(2, Int#(32)) _S16i25 = min_max(pack(s15[mod*i+25]) , pack(s15[mod*i+25+mod/2]));
			 Vector#(2, Int#(32)) _S16i26 = min_max(pack(s15[mod*i+26]) , pack(s15[mod*i+26+mod/2]));
			 Vector#(2, Int#(32)) _S16i27 = min_max(pack(s15[mod*i+27]) , pack(s15[mod*i+27+mod/2]));
			 Vector#(2, Int#(32)) _S16i28 = min_max(pack(s15[mod*i+28]) , pack(s15[mod*i+28+mod/2]));
			 Vector#(2, Int#(32)) _S16i29 = min_max(pack(s15[mod*i+29]) , pack(s15[mod*i+29+mod/2]));
			 Vector#(2, Int#(32)) _S16i30 = min_max(pack(s15[mod*i+30]) , pack(s15[mod*i+30+mod/2]));
			 Vector#(2, Int#(32)) _S16i31 = min_max(pack(s15[mod*i+31]) , pack(s15[mod*i+31+mod/2]));
		if ((i/1)%2 == 0) begin
			s16[mod*i+0] <= _S16i0[0];
			s16[mod*i+0+mod/2] <= _S16i0[1];
			s16[mod*i+1] <= _S16i1[0];
			s16[mod*i+1+mod/2] <= _S16i1[1];
			s16[mod*i+2] <= _S16i2[0];
			s16[mod*i+2+mod/2] <= _S16i2[1];
			s16[mod*i+3] <= _S16i3[0];
			s16[mod*i+3+mod/2] <= _S16i3[1];
			s16[mod*i+4] <= _S16i4[0];
			s16[mod*i+4+mod/2] <= _S16i4[1];
			s16[mod*i+5] <= _S16i5[0];
			s16[mod*i+5+mod/2] <= _S16i5[1];
			s16[mod*i+6] <= _S16i6[0];
			s16[mod*i+6+mod/2] <= _S16i6[1];
			s16[mod*i+7] <= _S16i7[0];
			s16[mod*i+7+mod/2] <= _S16i7[1];
			s16[mod*i+8] <= _S16i8[0];
			s16[mod*i+8+mod/2] <= _S16i8[1];
			s16[mod*i+9] <= _S16i9[0];
			s16[mod*i+9+mod/2] <= _S16i9[1];
			s16[mod*i+10] <= _S16i10[0];
			s16[mod*i+10+mod/2] <= _S16i10[1];
			s16[mod*i+11] <= _S16i11[0];
			s16[mod*i+11+mod/2] <= _S16i11[1];
			s16[mod*i+12] <= _S16i12[0];
			s16[mod*i+12+mod/2] <= _S16i12[1];
			s16[mod*i+13] <= _S16i13[0];
			s16[mod*i+13+mod/2] <= _S16i13[1];
			s16[mod*i+14] <= _S16i14[0];
			s16[mod*i+14+mod/2] <= _S16i14[1];
			s16[mod*i+15] <= _S16i15[0];
			s16[mod*i+15+mod/2] <= _S16i15[1];
			s16[mod*i+16] <= _S16i16[0];
			s16[mod*i+16+mod/2] <= _S16i16[1];
			s16[mod*i+17] <= _S16i17[0];
			s16[mod*i+17+mod/2] <= _S16i17[1];
			s16[mod*i+18] <= _S16i18[0];
			s16[mod*i+18+mod/2] <= _S16i18[1];
			s16[mod*i+19] <= _S16i19[0];
			s16[mod*i+19+mod/2] <= _S16i19[1];
			s16[mod*i+20] <= _S16i20[0];
			s16[mod*i+20+mod/2] <= _S16i20[1];
			s16[mod*i+21] <= _S16i21[0];
			s16[mod*i+21+mod/2] <= _S16i21[1];
			s16[mod*i+22] <= _S16i22[0];
			s16[mod*i+22+mod/2] <= _S16i22[1];
			s16[mod*i+23] <= _S16i23[0];
			s16[mod*i+23+mod/2] <= _S16i23[1];
			s16[mod*i+24] <= _S16i24[0];
			s16[mod*i+24+mod/2] <= _S16i24[1];
			s16[mod*i+25] <= _S16i25[0];
			s16[mod*i+25+mod/2] <= _S16i25[1];
			s16[mod*i+26] <= _S16i26[0];
			s16[mod*i+26+mod/2] <= _S16i26[1];
			s16[mod*i+27] <= _S16i27[0];
			s16[mod*i+27+mod/2] <= _S16i27[1];
			s16[mod*i+28] <= _S16i28[0];
			s16[mod*i+28+mod/2] <= _S16i28[1];
			s16[mod*i+29] <= _S16i29[0];
			s16[mod*i+29+mod/2] <= _S16i29[1];
			s16[mod*i+30] <= _S16i30[0];
			s16[mod*i+30+mod/2] <= _S16i30[1];
			s16[mod*i+31] <= _S16i31[0];
			s16[mod*i+31+mod/2] <= _S16i31[1];
		end
		else begin
			s16[mod*i+0] <= _S16i0[1];
			s16[mod*i+0+mod/2] <= _S16i0[0];
			s16[mod*i+1] <= _S16i1[1];
			s16[mod*i+1+mod/2] <= _S16i1[0];
			s16[mod*i+2] <= _S16i2[1];
			s16[mod*i+2+mod/2] <= _S16i2[0];
			s16[mod*i+3] <= _S16i3[1];
			s16[mod*i+3+mod/2] <= _S16i3[0];
			s16[mod*i+4] <= _S16i4[1];
			s16[mod*i+4+mod/2] <= _S16i4[0];
			s16[mod*i+5] <= _S16i5[1];
			s16[mod*i+5+mod/2] <= _S16i5[0];
			s16[mod*i+6] <= _S16i6[1];
			s16[mod*i+6+mod/2] <= _S16i6[0];
			s16[mod*i+7] <= _S16i7[1];
			s16[mod*i+7+mod/2] <= _S16i7[0];
			s16[mod*i+8] <= _S16i8[1];
			s16[mod*i+8+mod/2] <= _S16i8[0];
			s16[mod*i+9] <= _S16i9[1];
			s16[mod*i+9+mod/2] <= _S16i9[0];
			s16[mod*i+10] <= _S16i10[1];
			s16[mod*i+10+mod/2] <= _S16i10[0];
			s16[mod*i+11] <= _S16i11[1];
			s16[mod*i+11+mod/2] <= _S16i11[0];
			s16[mod*i+12] <= _S16i12[1];
			s16[mod*i+12+mod/2] <= _S16i12[0];
			s16[mod*i+13] <= _S16i13[1];
			s16[mod*i+13+mod/2] <= _S16i13[0];
			s16[mod*i+14] <= _S16i14[1];
			s16[mod*i+14+mod/2] <= _S16i14[0];
			s16[mod*i+15] <= _S16i15[1];
			s16[mod*i+15+mod/2] <= _S16i15[0];
			s16[mod*i+16] <= _S16i16[1];
			s16[mod*i+16+mod/2] <= _S16i16[0];
			s16[mod*i+17] <= _S16i17[1];
			s16[mod*i+17+mod/2] <= _S16i17[0];
			s16[mod*i+18] <= _S16i18[1];
			s16[mod*i+18+mod/2] <= _S16i18[0];
			s16[mod*i+19] <= _S16i19[1];
			s16[mod*i+19+mod/2] <= _S16i19[0];
			s16[mod*i+20] <= _S16i20[1];
			s16[mod*i+20+mod/2] <= _S16i20[0];
			s16[mod*i+21] <= _S16i21[1];
			s16[mod*i+21+mod/2] <= _S16i21[0];
			s16[mod*i+22] <= _S16i22[1];
			s16[mod*i+22+mod/2] <= _S16i22[0];
			s16[mod*i+23] <= _S16i23[1];
			s16[mod*i+23+mod/2] <= _S16i23[0];
			s16[mod*i+24] <= _S16i24[1];
			s16[mod*i+24+mod/2] <= _S16i24[0];
			s16[mod*i+25] <= _S16i25[1];
			s16[mod*i+25+mod/2] <= _S16i25[0];
			s16[mod*i+26] <= _S16i26[1];
			s16[mod*i+26+mod/2] <= _S16i26[0];
			s16[mod*i+27] <= _S16i27[1];
			s16[mod*i+27+mod/2] <= _S16i27[0];
			s16[mod*i+28] <= _S16i28[1];
			s16[mod*i+28+mod/2] <= _S16i28[0];
			s16[mod*i+29] <= _S16i29[1];
			s16[mod*i+29+mod/2] <= _S16i29[0];
			s16[mod*i+30] <= _S16i30[1];
			s16[mod*i+30+mod/2] <= _S16i30[0];
			s16[mod*i+31] <= _S16i31[1];
			s16[mod*i+31+mod/2] <= _S16i31[0];
		end
	end
	p16.enq(1);
endrule
rule _Q55;
	p16.deq;
	let mod = 32;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S17i0 = min_max(pack(s16[mod*i+0]) , pack(s16[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S17i1 = min_max(pack(s16[mod*i+1]) , pack(s16[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S17i2 = min_max(pack(s16[mod*i+2]) , pack(s16[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S17i3 = min_max(pack(s16[mod*i+3]) , pack(s16[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S17i4 = min_max(pack(s16[mod*i+4]) , pack(s16[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S17i5 = min_max(pack(s16[mod*i+5]) , pack(s16[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S17i6 = min_max(pack(s16[mod*i+6]) , pack(s16[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S17i7 = min_max(pack(s16[mod*i+7]) , pack(s16[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S17i8 = min_max(pack(s16[mod*i+8]) , pack(s16[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S17i9 = min_max(pack(s16[mod*i+9]) , pack(s16[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S17i10 = min_max(pack(s16[mod*i+10]) , pack(s16[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S17i11 = min_max(pack(s16[mod*i+11]) , pack(s16[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S17i12 = min_max(pack(s16[mod*i+12]) , pack(s16[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S17i13 = min_max(pack(s16[mod*i+13]) , pack(s16[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S17i14 = min_max(pack(s16[mod*i+14]) , pack(s16[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S17i15 = min_max(pack(s16[mod*i+15]) , pack(s16[mod*i+15+mod/2]));
		if ((i/2)%2 == 0) begin
			s17[mod*i+0] <= _S17i0[0];
			s17[mod*i+0+mod/2] <= _S17i0[1];
			s17[mod*i+1] <= _S17i1[0];
			s17[mod*i+1+mod/2] <= _S17i1[1];
			s17[mod*i+2] <= _S17i2[0];
			s17[mod*i+2+mod/2] <= _S17i2[1];
			s17[mod*i+3] <= _S17i3[0];
			s17[mod*i+3+mod/2] <= _S17i3[1];
			s17[mod*i+4] <= _S17i4[0];
			s17[mod*i+4+mod/2] <= _S17i4[1];
			s17[mod*i+5] <= _S17i5[0];
			s17[mod*i+5+mod/2] <= _S17i5[1];
			s17[mod*i+6] <= _S17i6[0];
			s17[mod*i+6+mod/2] <= _S17i6[1];
			s17[mod*i+7] <= _S17i7[0];
			s17[mod*i+7+mod/2] <= _S17i7[1];
			s17[mod*i+8] <= _S17i8[0];
			s17[mod*i+8+mod/2] <= _S17i8[1];
			s17[mod*i+9] <= _S17i9[0];
			s17[mod*i+9+mod/2] <= _S17i9[1];
			s17[mod*i+10] <= _S17i10[0];
			s17[mod*i+10+mod/2] <= _S17i10[1];
			s17[mod*i+11] <= _S17i11[0];
			s17[mod*i+11+mod/2] <= _S17i11[1];
			s17[mod*i+12] <= _S17i12[0];
			s17[mod*i+12+mod/2] <= _S17i12[1];
			s17[mod*i+13] <= _S17i13[0];
			s17[mod*i+13+mod/2] <= _S17i13[1];
			s17[mod*i+14] <= _S17i14[0];
			s17[mod*i+14+mod/2] <= _S17i14[1];
			s17[mod*i+15] <= _S17i15[0];
			s17[mod*i+15+mod/2] <= _S17i15[1];
		end
		else begin
			s17[mod*i+0] <= _S17i0[1];
			s17[mod*i+0+mod/2] <= _S17i0[0];
			s17[mod*i+1] <= _S17i1[1];
			s17[mod*i+1+mod/2] <= _S17i1[0];
			s17[mod*i+2] <= _S17i2[1];
			s17[mod*i+2+mod/2] <= _S17i2[0];
			s17[mod*i+3] <= _S17i3[1];
			s17[mod*i+3+mod/2] <= _S17i3[0];
			s17[mod*i+4] <= _S17i4[1];
			s17[mod*i+4+mod/2] <= _S17i4[0];
			s17[mod*i+5] <= _S17i5[1];
			s17[mod*i+5+mod/2] <= _S17i5[0];
			s17[mod*i+6] <= _S17i6[1];
			s17[mod*i+6+mod/2] <= _S17i6[0];
			s17[mod*i+7] <= _S17i7[1];
			s17[mod*i+7+mod/2] <= _S17i7[0];
			s17[mod*i+8] <= _S17i8[1];
			s17[mod*i+8+mod/2] <= _S17i8[0];
			s17[mod*i+9] <= _S17i9[1];
			s17[mod*i+9+mod/2] <= _S17i9[0];
			s17[mod*i+10] <= _S17i10[1];
			s17[mod*i+10+mod/2] <= _S17i10[0];
			s17[mod*i+11] <= _S17i11[1];
			s17[mod*i+11+mod/2] <= _S17i11[0];
			s17[mod*i+12] <= _S17i12[1];
			s17[mod*i+12+mod/2] <= _S17i12[0];
			s17[mod*i+13] <= _S17i13[1];
			s17[mod*i+13+mod/2] <= _S17i13[0];
			s17[mod*i+14] <= _S17i14[1];
			s17[mod*i+14+mod/2] <= _S17i14[0];
			s17[mod*i+15] <= _S17i15[1];
			s17[mod*i+15+mod/2] <= _S17i15[0];
		end
	end
	p17.enq(1);
endrule
rule _Q54;
	p17.deq;
	let mod = 16;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S18i0 = min_max(pack(s17[mod*i+0]) , pack(s17[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S18i1 = min_max(pack(s17[mod*i+1]) , pack(s17[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S18i2 = min_max(pack(s17[mod*i+2]) , pack(s17[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S18i3 = min_max(pack(s17[mod*i+3]) , pack(s17[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S18i4 = min_max(pack(s17[mod*i+4]) , pack(s17[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S18i5 = min_max(pack(s17[mod*i+5]) , pack(s17[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S18i6 = min_max(pack(s17[mod*i+6]) , pack(s17[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S18i7 = min_max(pack(s17[mod*i+7]) , pack(s17[mod*i+7+mod/2]));
		if ((i/4)%2 == 0) begin
			s18[mod*i+0] <= _S18i0[0];
			s18[mod*i+0+mod/2] <= _S18i0[1];
			s18[mod*i+1] <= _S18i1[0];
			s18[mod*i+1+mod/2] <= _S18i1[1];
			s18[mod*i+2] <= _S18i2[0];
			s18[mod*i+2+mod/2] <= _S18i2[1];
			s18[mod*i+3] <= _S18i3[0];
			s18[mod*i+3+mod/2] <= _S18i3[1];
			s18[mod*i+4] <= _S18i4[0];
			s18[mod*i+4+mod/2] <= _S18i4[1];
			s18[mod*i+5] <= _S18i5[0];
			s18[mod*i+5+mod/2] <= _S18i5[1];
			s18[mod*i+6] <= _S18i6[0];
			s18[mod*i+6+mod/2] <= _S18i6[1];
			s18[mod*i+7] <= _S18i7[0];
			s18[mod*i+7+mod/2] <= _S18i7[1];
		end
		else begin
			s18[mod*i+0] <= _S18i0[1];
			s18[mod*i+0+mod/2] <= _S18i0[0];
			s18[mod*i+1] <= _S18i1[1];
			s18[mod*i+1+mod/2] <= _S18i1[0];
			s18[mod*i+2] <= _S18i2[1];
			s18[mod*i+2+mod/2] <= _S18i2[0];
			s18[mod*i+3] <= _S18i3[1];
			s18[mod*i+3+mod/2] <= _S18i3[0];
			s18[mod*i+4] <= _S18i4[1];
			s18[mod*i+4+mod/2] <= _S18i4[0];
			s18[mod*i+5] <= _S18i5[1];
			s18[mod*i+5+mod/2] <= _S18i5[0];
			s18[mod*i+6] <= _S18i6[1];
			s18[mod*i+6+mod/2] <= _S18i6[0];
			s18[mod*i+7] <= _S18i7[1];
			s18[mod*i+7+mod/2] <= _S18i7[0];
		end
	end
	p18.enq(1);
endrule
rule _Q53;
	p18.deq;
	let mod = 8;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S19i0 = min_max(pack(s18[mod*i+0]) , pack(s18[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S19i1 = min_max(pack(s18[mod*i+1]) , pack(s18[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S19i2 = min_max(pack(s18[mod*i+2]) , pack(s18[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S19i3 = min_max(pack(s18[mod*i+3]) , pack(s18[mod*i+3+mod/2]));
		if ((i/8)%2 == 0) begin
			s19[mod*i+0] <= _S19i0[0];
			s19[mod*i+0+mod/2] <= _S19i0[1];
			s19[mod*i+1] <= _S19i1[0];
			s19[mod*i+1+mod/2] <= _S19i1[1];
			s19[mod*i+2] <= _S19i2[0];
			s19[mod*i+2+mod/2] <= _S19i2[1];
			s19[mod*i+3] <= _S19i3[0];
			s19[mod*i+3+mod/2] <= _S19i3[1];
		end
		else begin
			s19[mod*i+0] <= _S19i0[1];
			s19[mod*i+0+mod/2] <= _S19i0[0];
			s19[mod*i+1] <= _S19i1[1];
			s19[mod*i+1+mod/2] <= _S19i1[0];
			s19[mod*i+2] <= _S19i2[1];
			s19[mod*i+2+mod/2] <= _S19i2[0];
			s19[mod*i+3] <= _S19i3[1];
			s19[mod*i+3+mod/2] <= _S19i3[0];
		end
	end
	p19.enq(1);
endrule
rule _Q52;
	p19.deq;
	let mod = 4;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S20i0 = min_max(pack(s19[mod*i+0]) , pack(s19[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S20i1 = min_max(pack(s19[mod*i+1]) , pack(s19[mod*i+1+mod/2]));
		if ((i/16)%2 == 0) begin
			s20[mod*i+0] <= _S20i0[0];
			s20[mod*i+0+mod/2] <= _S20i0[1];
			s20[mod*i+1] <= _S20i1[0];
			s20[mod*i+1+mod/2] <= _S20i1[1];
		end
		else begin
			s20[mod*i+0] <= _S20i0[1];
			s20[mod*i+0+mod/2] <= _S20i0[0];
			s20[mod*i+1] <= _S20i1[1];
			s20[mod*i+1+mod/2] <= _S20i1[0];
		end
	end
	p20.enq(1);
endrule
rule _Q51;
	p20.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S21i0 = min_max(pack(s20[mod*i+0]) , pack(s20[mod*i+0+mod/2]));
		if ((i/32)%2 == 0) begin
			s21[mod*i+0] <= _S21i0[0];
			s21[mod*i+0+mod/2] <= _S21i0[1];
		end
		else begin
			s21[mod*i+0] <= _S21i0[1];
			s21[mod*i+0+mod/2] <= _S21i0[0];
		end
	end
	p21.enq(1);
endrule
rule _Q67;
	p21.deq;
	let mod = 128;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S22i0 = min_max(pack(s21[mod*i+0]) , pack(s21[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S22i1 = min_max(pack(s21[mod*i+1]) , pack(s21[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S22i2 = min_max(pack(s21[mod*i+2]) , pack(s21[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S22i3 = min_max(pack(s21[mod*i+3]) , pack(s21[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S22i4 = min_max(pack(s21[mod*i+4]) , pack(s21[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S22i5 = min_max(pack(s21[mod*i+5]) , pack(s21[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S22i6 = min_max(pack(s21[mod*i+6]) , pack(s21[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S22i7 = min_max(pack(s21[mod*i+7]) , pack(s21[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S22i8 = min_max(pack(s21[mod*i+8]) , pack(s21[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S22i9 = min_max(pack(s21[mod*i+9]) , pack(s21[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S22i10 = min_max(pack(s21[mod*i+10]) , pack(s21[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S22i11 = min_max(pack(s21[mod*i+11]) , pack(s21[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S22i12 = min_max(pack(s21[mod*i+12]) , pack(s21[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S22i13 = min_max(pack(s21[mod*i+13]) , pack(s21[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S22i14 = min_max(pack(s21[mod*i+14]) , pack(s21[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S22i15 = min_max(pack(s21[mod*i+15]) , pack(s21[mod*i+15+mod/2]));
			 Vector#(2, Int#(32)) _S22i16 = min_max(pack(s21[mod*i+16]) , pack(s21[mod*i+16+mod/2]));
			 Vector#(2, Int#(32)) _S22i17 = min_max(pack(s21[mod*i+17]) , pack(s21[mod*i+17+mod/2]));
			 Vector#(2, Int#(32)) _S22i18 = min_max(pack(s21[mod*i+18]) , pack(s21[mod*i+18+mod/2]));
			 Vector#(2, Int#(32)) _S22i19 = min_max(pack(s21[mod*i+19]) , pack(s21[mod*i+19+mod/2]));
			 Vector#(2, Int#(32)) _S22i20 = min_max(pack(s21[mod*i+20]) , pack(s21[mod*i+20+mod/2]));
			 Vector#(2, Int#(32)) _S22i21 = min_max(pack(s21[mod*i+21]) , pack(s21[mod*i+21+mod/2]));
			 Vector#(2, Int#(32)) _S22i22 = min_max(pack(s21[mod*i+22]) , pack(s21[mod*i+22+mod/2]));
			 Vector#(2, Int#(32)) _S22i23 = min_max(pack(s21[mod*i+23]) , pack(s21[mod*i+23+mod/2]));
			 Vector#(2, Int#(32)) _S22i24 = min_max(pack(s21[mod*i+24]) , pack(s21[mod*i+24+mod/2]));
			 Vector#(2, Int#(32)) _S22i25 = min_max(pack(s21[mod*i+25]) , pack(s21[mod*i+25+mod/2]));
			 Vector#(2, Int#(32)) _S22i26 = min_max(pack(s21[mod*i+26]) , pack(s21[mod*i+26+mod/2]));
			 Vector#(2, Int#(32)) _S22i27 = min_max(pack(s21[mod*i+27]) , pack(s21[mod*i+27+mod/2]));
			 Vector#(2, Int#(32)) _S22i28 = min_max(pack(s21[mod*i+28]) , pack(s21[mod*i+28+mod/2]));
			 Vector#(2, Int#(32)) _S22i29 = min_max(pack(s21[mod*i+29]) , pack(s21[mod*i+29+mod/2]));
			 Vector#(2, Int#(32)) _S22i30 = min_max(pack(s21[mod*i+30]) , pack(s21[mod*i+30+mod/2]));
			 Vector#(2, Int#(32)) _S22i31 = min_max(pack(s21[mod*i+31]) , pack(s21[mod*i+31+mod/2]));
			 Vector#(2, Int#(32)) _S22i32 = min_max(pack(s21[mod*i+32]) , pack(s21[mod*i+32+mod/2]));
			 Vector#(2, Int#(32)) _S22i33 = min_max(pack(s21[mod*i+33]) , pack(s21[mod*i+33+mod/2]));
			 Vector#(2, Int#(32)) _S22i34 = min_max(pack(s21[mod*i+34]) , pack(s21[mod*i+34+mod/2]));
			 Vector#(2, Int#(32)) _S22i35 = min_max(pack(s21[mod*i+35]) , pack(s21[mod*i+35+mod/2]));
			 Vector#(2, Int#(32)) _S22i36 = min_max(pack(s21[mod*i+36]) , pack(s21[mod*i+36+mod/2]));
			 Vector#(2, Int#(32)) _S22i37 = min_max(pack(s21[mod*i+37]) , pack(s21[mod*i+37+mod/2]));
			 Vector#(2, Int#(32)) _S22i38 = min_max(pack(s21[mod*i+38]) , pack(s21[mod*i+38+mod/2]));
			 Vector#(2, Int#(32)) _S22i39 = min_max(pack(s21[mod*i+39]) , pack(s21[mod*i+39+mod/2]));
			 Vector#(2, Int#(32)) _S22i40 = min_max(pack(s21[mod*i+40]) , pack(s21[mod*i+40+mod/2]));
			 Vector#(2, Int#(32)) _S22i41 = min_max(pack(s21[mod*i+41]) , pack(s21[mod*i+41+mod/2]));
			 Vector#(2, Int#(32)) _S22i42 = min_max(pack(s21[mod*i+42]) , pack(s21[mod*i+42+mod/2]));
			 Vector#(2, Int#(32)) _S22i43 = min_max(pack(s21[mod*i+43]) , pack(s21[mod*i+43+mod/2]));
			 Vector#(2, Int#(32)) _S22i44 = min_max(pack(s21[mod*i+44]) , pack(s21[mod*i+44+mod/2]));
			 Vector#(2, Int#(32)) _S22i45 = min_max(pack(s21[mod*i+45]) , pack(s21[mod*i+45+mod/2]));
			 Vector#(2, Int#(32)) _S22i46 = min_max(pack(s21[mod*i+46]) , pack(s21[mod*i+46+mod/2]));
			 Vector#(2, Int#(32)) _S22i47 = min_max(pack(s21[mod*i+47]) , pack(s21[mod*i+47+mod/2]));
			 Vector#(2, Int#(32)) _S22i48 = min_max(pack(s21[mod*i+48]) , pack(s21[mod*i+48+mod/2]));
			 Vector#(2, Int#(32)) _S22i49 = min_max(pack(s21[mod*i+49]) , pack(s21[mod*i+49+mod/2]));
			 Vector#(2, Int#(32)) _S22i50 = min_max(pack(s21[mod*i+50]) , pack(s21[mod*i+50+mod/2]));
			 Vector#(2, Int#(32)) _S22i51 = min_max(pack(s21[mod*i+51]) , pack(s21[mod*i+51+mod/2]));
			 Vector#(2, Int#(32)) _S22i52 = min_max(pack(s21[mod*i+52]) , pack(s21[mod*i+52+mod/2]));
			 Vector#(2, Int#(32)) _S22i53 = min_max(pack(s21[mod*i+53]) , pack(s21[mod*i+53+mod/2]));
			 Vector#(2, Int#(32)) _S22i54 = min_max(pack(s21[mod*i+54]) , pack(s21[mod*i+54+mod/2]));
			 Vector#(2, Int#(32)) _S22i55 = min_max(pack(s21[mod*i+55]) , pack(s21[mod*i+55+mod/2]));
			 Vector#(2, Int#(32)) _S22i56 = min_max(pack(s21[mod*i+56]) , pack(s21[mod*i+56+mod/2]));
			 Vector#(2, Int#(32)) _S22i57 = min_max(pack(s21[mod*i+57]) , pack(s21[mod*i+57+mod/2]));
			 Vector#(2, Int#(32)) _S22i58 = min_max(pack(s21[mod*i+58]) , pack(s21[mod*i+58+mod/2]));
			 Vector#(2, Int#(32)) _S22i59 = min_max(pack(s21[mod*i+59]) , pack(s21[mod*i+59+mod/2]));
			 Vector#(2, Int#(32)) _S22i60 = min_max(pack(s21[mod*i+60]) , pack(s21[mod*i+60+mod/2]));
			 Vector#(2, Int#(32)) _S22i61 = min_max(pack(s21[mod*i+61]) , pack(s21[mod*i+61+mod/2]));
			 Vector#(2, Int#(32)) _S22i62 = min_max(pack(s21[mod*i+62]) , pack(s21[mod*i+62+mod/2]));
			 Vector#(2, Int#(32)) _S22i63 = min_max(pack(s21[mod*i+63]) , pack(s21[mod*i+63+mod/2]));
		if ((i/1)%2 == 0) begin
			s22[mod*i+0] <= _S22i0[0];
			s22[mod*i+0+mod/2] <= _S22i0[1];
			s22[mod*i+1] <= _S22i1[0];
			s22[mod*i+1+mod/2] <= _S22i1[1];
			s22[mod*i+2] <= _S22i2[0];
			s22[mod*i+2+mod/2] <= _S22i2[1];
			s22[mod*i+3] <= _S22i3[0];
			s22[mod*i+3+mod/2] <= _S22i3[1];
			s22[mod*i+4] <= _S22i4[0];
			s22[mod*i+4+mod/2] <= _S22i4[1];
			s22[mod*i+5] <= _S22i5[0];
			s22[mod*i+5+mod/2] <= _S22i5[1];
			s22[mod*i+6] <= _S22i6[0];
			s22[mod*i+6+mod/2] <= _S22i6[1];
			s22[mod*i+7] <= _S22i7[0];
			s22[mod*i+7+mod/2] <= _S22i7[1];
			s22[mod*i+8] <= _S22i8[0];
			s22[mod*i+8+mod/2] <= _S22i8[1];
			s22[mod*i+9] <= _S22i9[0];
			s22[mod*i+9+mod/2] <= _S22i9[1];
			s22[mod*i+10] <= _S22i10[0];
			s22[mod*i+10+mod/2] <= _S22i10[1];
			s22[mod*i+11] <= _S22i11[0];
			s22[mod*i+11+mod/2] <= _S22i11[1];
			s22[mod*i+12] <= _S22i12[0];
			s22[mod*i+12+mod/2] <= _S22i12[1];
			s22[mod*i+13] <= _S22i13[0];
			s22[mod*i+13+mod/2] <= _S22i13[1];
			s22[mod*i+14] <= _S22i14[0];
			s22[mod*i+14+mod/2] <= _S22i14[1];
			s22[mod*i+15] <= _S22i15[0];
			s22[mod*i+15+mod/2] <= _S22i15[1];
			s22[mod*i+16] <= _S22i16[0];
			s22[mod*i+16+mod/2] <= _S22i16[1];
			s22[mod*i+17] <= _S22i17[0];
			s22[mod*i+17+mod/2] <= _S22i17[1];
			s22[mod*i+18] <= _S22i18[0];
			s22[mod*i+18+mod/2] <= _S22i18[1];
			s22[mod*i+19] <= _S22i19[0];
			s22[mod*i+19+mod/2] <= _S22i19[1];
			s22[mod*i+20] <= _S22i20[0];
			s22[mod*i+20+mod/2] <= _S22i20[1];
			s22[mod*i+21] <= _S22i21[0];
			s22[mod*i+21+mod/2] <= _S22i21[1];
			s22[mod*i+22] <= _S22i22[0];
			s22[mod*i+22+mod/2] <= _S22i22[1];
			s22[mod*i+23] <= _S22i23[0];
			s22[mod*i+23+mod/2] <= _S22i23[1];
			s22[mod*i+24] <= _S22i24[0];
			s22[mod*i+24+mod/2] <= _S22i24[1];
			s22[mod*i+25] <= _S22i25[0];
			s22[mod*i+25+mod/2] <= _S22i25[1];
			s22[mod*i+26] <= _S22i26[0];
			s22[mod*i+26+mod/2] <= _S22i26[1];
			s22[mod*i+27] <= _S22i27[0];
			s22[mod*i+27+mod/2] <= _S22i27[1];
			s22[mod*i+28] <= _S22i28[0];
			s22[mod*i+28+mod/2] <= _S22i28[1];
			s22[mod*i+29] <= _S22i29[0];
			s22[mod*i+29+mod/2] <= _S22i29[1];
			s22[mod*i+30] <= _S22i30[0];
			s22[mod*i+30+mod/2] <= _S22i30[1];
			s22[mod*i+31] <= _S22i31[0];
			s22[mod*i+31+mod/2] <= _S22i31[1];
			s22[mod*i+32] <= _S22i32[0];
			s22[mod*i+32+mod/2] <= _S22i32[1];
			s22[mod*i+33] <= _S22i33[0];
			s22[mod*i+33+mod/2] <= _S22i33[1];
			s22[mod*i+34] <= _S22i34[0];
			s22[mod*i+34+mod/2] <= _S22i34[1];
			s22[mod*i+35] <= _S22i35[0];
			s22[mod*i+35+mod/2] <= _S22i35[1];
			s22[mod*i+36] <= _S22i36[0];
			s22[mod*i+36+mod/2] <= _S22i36[1];
			s22[mod*i+37] <= _S22i37[0];
			s22[mod*i+37+mod/2] <= _S22i37[1];
			s22[mod*i+38] <= _S22i38[0];
			s22[mod*i+38+mod/2] <= _S22i38[1];
			s22[mod*i+39] <= _S22i39[0];
			s22[mod*i+39+mod/2] <= _S22i39[1];
			s22[mod*i+40] <= _S22i40[0];
			s22[mod*i+40+mod/2] <= _S22i40[1];
			s22[mod*i+41] <= _S22i41[0];
			s22[mod*i+41+mod/2] <= _S22i41[1];
			s22[mod*i+42] <= _S22i42[0];
			s22[mod*i+42+mod/2] <= _S22i42[1];
			s22[mod*i+43] <= _S22i43[0];
			s22[mod*i+43+mod/2] <= _S22i43[1];
			s22[mod*i+44] <= _S22i44[0];
			s22[mod*i+44+mod/2] <= _S22i44[1];
			s22[mod*i+45] <= _S22i45[0];
			s22[mod*i+45+mod/2] <= _S22i45[1];
			s22[mod*i+46] <= _S22i46[0];
			s22[mod*i+46+mod/2] <= _S22i46[1];
			s22[mod*i+47] <= _S22i47[0];
			s22[mod*i+47+mod/2] <= _S22i47[1];
			s22[mod*i+48] <= _S22i48[0];
			s22[mod*i+48+mod/2] <= _S22i48[1];
			s22[mod*i+49] <= _S22i49[0];
			s22[mod*i+49+mod/2] <= _S22i49[1];
			s22[mod*i+50] <= _S22i50[0];
			s22[mod*i+50+mod/2] <= _S22i50[1];
			s22[mod*i+51] <= _S22i51[0];
			s22[mod*i+51+mod/2] <= _S22i51[1];
			s22[mod*i+52] <= _S22i52[0];
			s22[mod*i+52+mod/2] <= _S22i52[1];
			s22[mod*i+53] <= _S22i53[0];
			s22[mod*i+53+mod/2] <= _S22i53[1];
			s22[mod*i+54] <= _S22i54[0];
			s22[mod*i+54+mod/2] <= _S22i54[1];
			s22[mod*i+55] <= _S22i55[0];
			s22[mod*i+55+mod/2] <= _S22i55[1];
			s22[mod*i+56] <= _S22i56[0];
			s22[mod*i+56+mod/2] <= _S22i56[1];
			s22[mod*i+57] <= _S22i57[0];
			s22[mod*i+57+mod/2] <= _S22i57[1];
			s22[mod*i+58] <= _S22i58[0];
			s22[mod*i+58+mod/2] <= _S22i58[1];
			s22[mod*i+59] <= _S22i59[0];
			s22[mod*i+59+mod/2] <= _S22i59[1];
			s22[mod*i+60] <= _S22i60[0];
			s22[mod*i+60+mod/2] <= _S22i60[1];
			s22[mod*i+61] <= _S22i61[0];
			s22[mod*i+61+mod/2] <= _S22i61[1];
			s22[mod*i+62] <= _S22i62[0];
			s22[mod*i+62+mod/2] <= _S22i62[1];
			s22[mod*i+63] <= _S22i63[0];
			s22[mod*i+63+mod/2] <= _S22i63[1];
		end
		else begin
			s22[mod*i+0] <= _S22i0[1];
			s22[mod*i+0+mod/2] <= _S22i0[0];
			s22[mod*i+1] <= _S22i1[1];
			s22[mod*i+1+mod/2] <= _S22i1[0];
			s22[mod*i+2] <= _S22i2[1];
			s22[mod*i+2+mod/2] <= _S22i2[0];
			s22[mod*i+3] <= _S22i3[1];
			s22[mod*i+3+mod/2] <= _S22i3[0];
			s22[mod*i+4] <= _S22i4[1];
			s22[mod*i+4+mod/2] <= _S22i4[0];
			s22[mod*i+5] <= _S22i5[1];
			s22[mod*i+5+mod/2] <= _S22i5[0];
			s22[mod*i+6] <= _S22i6[1];
			s22[mod*i+6+mod/2] <= _S22i6[0];
			s22[mod*i+7] <= _S22i7[1];
			s22[mod*i+7+mod/2] <= _S22i7[0];
			s22[mod*i+8] <= _S22i8[1];
			s22[mod*i+8+mod/2] <= _S22i8[0];
			s22[mod*i+9] <= _S22i9[1];
			s22[mod*i+9+mod/2] <= _S22i9[0];
			s22[mod*i+10] <= _S22i10[1];
			s22[mod*i+10+mod/2] <= _S22i10[0];
			s22[mod*i+11] <= _S22i11[1];
			s22[mod*i+11+mod/2] <= _S22i11[0];
			s22[mod*i+12] <= _S22i12[1];
			s22[mod*i+12+mod/2] <= _S22i12[0];
			s22[mod*i+13] <= _S22i13[1];
			s22[mod*i+13+mod/2] <= _S22i13[0];
			s22[mod*i+14] <= _S22i14[1];
			s22[mod*i+14+mod/2] <= _S22i14[0];
			s22[mod*i+15] <= _S22i15[1];
			s22[mod*i+15+mod/2] <= _S22i15[0];
			s22[mod*i+16] <= _S22i16[1];
			s22[mod*i+16+mod/2] <= _S22i16[0];
			s22[mod*i+17] <= _S22i17[1];
			s22[mod*i+17+mod/2] <= _S22i17[0];
			s22[mod*i+18] <= _S22i18[1];
			s22[mod*i+18+mod/2] <= _S22i18[0];
			s22[mod*i+19] <= _S22i19[1];
			s22[mod*i+19+mod/2] <= _S22i19[0];
			s22[mod*i+20] <= _S22i20[1];
			s22[mod*i+20+mod/2] <= _S22i20[0];
			s22[mod*i+21] <= _S22i21[1];
			s22[mod*i+21+mod/2] <= _S22i21[0];
			s22[mod*i+22] <= _S22i22[1];
			s22[mod*i+22+mod/2] <= _S22i22[0];
			s22[mod*i+23] <= _S22i23[1];
			s22[mod*i+23+mod/2] <= _S22i23[0];
			s22[mod*i+24] <= _S22i24[1];
			s22[mod*i+24+mod/2] <= _S22i24[0];
			s22[mod*i+25] <= _S22i25[1];
			s22[mod*i+25+mod/2] <= _S22i25[0];
			s22[mod*i+26] <= _S22i26[1];
			s22[mod*i+26+mod/2] <= _S22i26[0];
			s22[mod*i+27] <= _S22i27[1];
			s22[mod*i+27+mod/2] <= _S22i27[0];
			s22[mod*i+28] <= _S22i28[1];
			s22[mod*i+28+mod/2] <= _S22i28[0];
			s22[mod*i+29] <= _S22i29[1];
			s22[mod*i+29+mod/2] <= _S22i29[0];
			s22[mod*i+30] <= _S22i30[1];
			s22[mod*i+30+mod/2] <= _S22i30[0];
			s22[mod*i+31] <= _S22i31[1];
			s22[mod*i+31+mod/2] <= _S22i31[0];
			s22[mod*i+32] <= _S22i32[1];
			s22[mod*i+32+mod/2] <= _S22i32[0];
			s22[mod*i+33] <= _S22i33[1];
			s22[mod*i+33+mod/2] <= _S22i33[0];
			s22[mod*i+34] <= _S22i34[1];
			s22[mod*i+34+mod/2] <= _S22i34[0];
			s22[mod*i+35] <= _S22i35[1];
			s22[mod*i+35+mod/2] <= _S22i35[0];
			s22[mod*i+36] <= _S22i36[1];
			s22[mod*i+36+mod/2] <= _S22i36[0];
			s22[mod*i+37] <= _S22i37[1];
			s22[mod*i+37+mod/2] <= _S22i37[0];
			s22[mod*i+38] <= _S22i38[1];
			s22[mod*i+38+mod/2] <= _S22i38[0];
			s22[mod*i+39] <= _S22i39[1];
			s22[mod*i+39+mod/2] <= _S22i39[0];
			s22[mod*i+40] <= _S22i40[1];
			s22[mod*i+40+mod/2] <= _S22i40[0];
			s22[mod*i+41] <= _S22i41[1];
			s22[mod*i+41+mod/2] <= _S22i41[0];
			s22[mod*i+42] <= _S22i42[1];
			s22[mod*i+42+mod/2] <= _S22i42[0];
			s22[mod*i+43] <= _S22i43[1];
			s22[mod*i+43+mod/2] <= _S22i43[0];
			s22[mod*i+44] <= _S22i44[1];
			s22[mod*i+44+mod/2] <= _S22i44[0];
			s22[mod*i+45] <= _S22i45[1];
			s22[mod*i+45+mod/2] <= _S22i45[0];
			s22[mod*i+46] <= _S22i46[1];
			s22[mod*i+46+mod/2] <= _S22i46[0];
			s22[mod*i+47] <= _S22i47[1];
			s22[mod*i+47+mod/2] <= _S22i47[0];
			s22[mod*i+48] <= _S22i48[1];
			s22[mod*i+48+mod/2] <= _S22i48[0];
			s22[mod*i+49] <= _S22i49[1];
			s22[mod*i+49+mod/2] <= _S22i49[0];
			s22[mod*i+50] <= _S22i50[1];
			s22[mod*i+50+mod/2] <= _S22i50[0];
			s22[mod*i+51] <= _S22i51[1];
			s22[mod*i+51+mod/2] <= _S22i51[0];
			s22[mod*i+52] <= _S22i52[1];
			s22[mod*i+52+mod/2] <= _S22i52[0];
			s22[mod*i+53] <= _S22i53[1];
			s22[mod*i+53+mod/2] <= _S22i53[0];
			s22[mod*i+54] <= _S22i54[1];
			s22[mod*i+54+mod/2] <= _S22i54[0];
			s22[mod*i+55] <= _S22i55[1];
			s22[mod*i+55+mod/2] <= _S22i55[0];
			s22[mod*i+56] <= _S22i56[1];
			s22[mod*i+56+mod/2] <= _S22i56[0];
			s22[mod*i+57] <= _S22i57[1];
			s22[mod*i+57+mod/2] <= _S22i57[0];
			s22[mod*i+58] <= _S22i58[1];
			s22[mod*i+58+mod/2] <= _S22i58[0];
			s22[mod*i+59] <= _S22i59[1];
			s22[mod*i+59+mod/2] <= _S22i59[0];
			s22[mod*i+60] <= _S22i60[1];
			s22[mod*i+60+mod/2] <= _S22i60[0];
			s22[mod*i+61] <= _S22i61[1];
			s22[mod*i+61+mod/2] <= _S22i61[0];
			s22[mod*i+62] <= _S22i62[1];
			s22[mod*i+62+mod/2] <= _S22i62[0];
			s22[mod*i+63] <= _S22i63[1];
			s22[mod*i+63+mod/2] <= _S22i63[0];
		end
	end
	p22.enq(1);
endrule
rule _Q66;
	p22.deq;
	let mod = 64;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S23i0 = min_max(pack(s22[mod*i+0]) , pack(s22[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S23i1 = min_max(pack(s22[mod*i+1]) , pack(s22[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S23i2 = min_max(pack(s22[mod*i+2]) , pack(s22[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S23i3 = min_max(pack(s22[mod*i+3]) , pack(s22[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S23i4 = min_max(pack(s22[mod*i+4]) , pack(s22[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S23i5 = min_max(pack(s22[mod*i+5]) , pack(s22[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S23i6 = min_max(pack(s22[mod*i+6]) , pack(s22[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S23i7 = min_max(pack(s22[mod*i+7]) , pack(s22[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S23i8 = min_max(pack(s22[mod*i+8]) , pack(s22[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S23i9 = min_max(pack(s22[mod*i+9]) , pack(s22[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S23i10 = min_max(pack(s22[mod*i+10]) , pack(s22[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S23i11 = min_max(pack(s22[mod*i+11]) , pack(s22[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S23i12 = min_max(pack(s22[mod*i+12]) , pack(s22[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S23i13 = min_max(pack(s22[mod*i+13]) , pack(s22[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S23i14 = min_max(pack(s22[mod*i+14]) , pack(s22[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S23i15 = min_max(pack(s22[mod*i+15]) , pack(s22[mod*i+15+mod/2]));
			 Vector#(2, Int#(32)) _S23i16 = min_max(pack(s22[mod*i+16]) , pack(s22[mod*i+16+mod/2]));
			 Vector#(2, Int#(32)) _S23i17 = min_max(pack(s22[mod*i+17]) , pack(s22[mod*i+17+mod/2]));
			 Vector#(2, Int#(32)) _S23i18 = min_max(pack(s22[mod*i+18]) , pack(s22[mod*i+18+mod/2]));
			 Vector#(2, Int#(32)) _S23i19 = min_max(pack(s22[mod*i+19]) , pack(s22[mod*i+19+mod/2]));
			 Vector#(2, Int#(32)) _S23i20 = min_max(pack(s22[mod*i+20]) , pack(s22[mod*i+20+mod/2]));
			 Vector#(2, Int#(32)) _S23i21 = min_max(pack(s22[mod*i+21]) , pack(s22[mod*i+21+mod/2]));
			 Vector#(2, Int#(32)) _S23i22 = min_max(pack(s22[mod*i+22]) , pack(s22[mod*i+22+mod/2]));
			 Vector#(2, Int#(32)) _S23i23 = min_max(pack(s22[mod*i+23]) , pack(s22[mod*i+23+mod/2]));
			 Vector#(2, Int#(32)) _S23i24 = min_max(pack(s22[mod*i+24]) , pack(s22[mod*i+24+mod/2]));
			 Vector#(2, Int#(32)) _S23i25 = min_max(pack(s22[mod*i+25]) , pack(s22[mod*i+25+mod/2]));
			 Vector#(2, Int#(32)) _S23i26 = min_max(pack(s22[mod*i+26]) , pack(s22[mod*i+26+mod/2]));
			 Vector#(2, Int#(32)) _S23i27 = min_max(pack(s22[mod*i+27]) , pack(s22[mod*i+27+mod/2]));
			 Vector#(2, Int#(32)) _S23i28 = min_max(pack(s22[mod*i+28]) , pack(s22[mod*i+28+mod/2]));
			 Vector#(2, Int#(32)) _S23i29 = min_max(pack(s22[mod*i+29]) , pack(s22[mod*i+29+mod/2]));
			 Vector#(2, Int#(32)) _S23i30 = min_max(pack(s22[mod*i+30]) , pack(s22[mod*i+30+mod/2]));
			 Vector#(2, Int#(32)) _S23i31 = min_max(pack(s22[mod*i+31]) , pack(s22[mod*i+31+mod/2]));
		if ((i/2)%2 == 0) begin
			s23[mod*i+0] <= _S23i0[0];
			s23[mod*i+0+mod/2] <= _S23i0[1];
			s23[mod*i+1] <= _S23i1[0];
			s23[mod*i+1+mod/2] <= _S23i1[1];
			s23[mod*i+2] <= _S23i2[0];
			s23[mod*i+2+mod/2] <= _S23i2[1];
			s23[mod*i+3] <= _S23i3[0];
			s23[mod*i+3+mod/2] <= _S23i3[1];
			s23[mod*i+4] <= _S23i4[0];
			s23[mod*i+4+mod/2] <= _S23i4[1];
			s23[mod*i+5] <= _S23i5[0];
			s23[mod*i+5+mod/2] <= _S23i5[1];
			s23[mod*i+6] <= _S23i6[0];
			s23[mod*i+6+mod/2] <= _S23i6[1];
			s23[mod*i+7] <= _S23i7[0];
			s23[mod*i+7+mod/2] <= _S23i7[1];
			s23[mod*i+8] <= _S23i8[0];
			s23[mod*i+8+mod/2] <= _S23i8[1];
			s23[mod*i+9] <= _S23i9[0];
			s23[mod*i+9+mod/2] <= _S23i9[1];
			s23[mod*i+10] <= _S23i10[0];
			s23[mod*i+10+mod/2] <= _S23i10[1];
			s23[mod*i+11] <= _S23i11[0];
			s23[mod*i+11+mod/2] <= _S23i11[1];
			s23[mod*i+12] <= _S23i12[0];
			s23[mod*i+12+mod/2] <= _S23i12[1];
			s23[mod*i+13] <= _S23i13[0];
			s23[mod*i+13+mod/2] <= _S23i13[1];
			s23[mod*i+14] <= _S23i14[0];
			s23[mod*i+14+mod/2] <= _S23i14[1];
			s23[mod*i+15] <= _S23i15[0];
			s23[mod*i+15+mod/2] <= _S23i15[1];
			s23[mod*i+16] <= _S23i16[0];
			s23[mod*i+16+mod/2] <= _S23i16[1];
			s23[mod*i+17] <= _S23i17[0];
			s23[mod*i+17+mod/2] <= _S23i17[1];
			s23[mod*i+18] <= _S23i18[0];
			s23[mod*i+18+mod/2] <= _S23i18[1];
			s23[mod*i+19] <= _S23i19[0];
			s23[mod*i+19+mod/2] <= _S23i19[1];
			s23[mod*i+20] <= _S23i20[0];
			s23[mod*i+20+mod/2] <= _S23i20[1];
			s23[mod*i+21] <= _S23i21[0];
			s23[mod*i+21+mod/2] <= _S23i21[1];
			s23[mod*i+22] <= _S23i22[0];
			s23[mod*i+22+mod/2] <= _S23i22[1];
			s23[mod*i+23] <= _S23i23[0];
			s23[mod*i+23+mod/2] <= _S23i23[1];
			s23[mod*i+24] <= _S23i24[0];
			s23[mod*i+24+mod/2] <= _S23i24[1];
			s23[mod*i+25] <= _S23i25[0];
			s23[mod*i+25+mod/2] <= _S23i25[1];
			s23[mod*i+26] <= _S23i26[0];
			s23[mod*i+26+mod/2] <= _S23i26[1];
			s23[mod*i+27] <= _S23i27[0];
			s23[mod*i+27+mod/2] <= _S23i27[1];
			s23[mod*i+28] <= _S23i28[0];
			s23[mod*i+28+mod/2] <= _S23i28[1];
			s23[mod*i+29] <= _S23i29[0];
			s23[mod*i+29+mod/2] <= _S23i29[1];
			s23[mod*i+30] <= _S23i30[0];
			s23[mod*i+30+mod/2] <= _S23i30[1];
			s23[mod*i+31] <= _S23i31[0];
			s23[mod*i+31+mod/2] <= _S23i31[1];
		end
		else begin
			s23[mod*i+0] <= _S23i0[1];
			s23[mod*i+0+mod/2] <= _S23i0[0];
			s23[mod*i+1] <= _S23i1[1];
			s23[mod*i+1+mod/2] <= _S23i1[0];
			s23[mod*i+2] <= _S23i2[1];
			s23[mod*i+2+mod/2] <= _S23i2[0];
			s23[mod*i+3] <= _S23i3[1];
			s23[mod*i+3+mod/2] <= _S23i3[0];
			s23[mod*i+4] <= _S23i4[1];
			s23[mod*i+4+mod/2] <= _S23i4[0];
			s23[mod*i+5] <= _S23i5[1];
			s23[mod*i+5+mod/2] <= _S23i5[0];
			s23[mod*i+6] <= _S23i6[1];
			s23[mod*i+6+mod/2] <= _S23i6[0];
			s23[mod*i+7] <= _S23i7[1];
			s23[mod*i+7+mod/2] <= _S23i7[0];
			s23[mod*i+8] <= _S23i8[1];
			s23[mod*i+8+mod/2] <= _S23i8[0];
			s23[mod*i+9] <= _S23i9[1];
			s23[mod*i+9+mod/2] <= _S23i9[0];
			s23[mod*i+10] <= _S23i10[1];
			s23[mod*i+10+mod/2] <= _S23i10[0];
			s23[mod*i+11] <= _S23i11[1];
			s23[mod*i+11+mod/2] <= _S23i11[0];
			s23[mod*i+12] <= _S23i12[1];
			s23[mod*i+12+mod/2] <= _S23i12[0];
			s23[mod*i+13] <= _S23i13[1];
			s23[mod*i+13+mod/2] <= _S23i13[0];
			s23[mod*i+14] <= _S23i14[1];
			s23[mod*i+14+mod/2] <= _S23i14[0];
			s23[mod*i+15] <= _S23i15[1];
			s23[mod*i+15+mod/2] <= _S23i15[0];
			s23[mod*i+16] <= _S23i16[1];
			s23[mod*i+16+mod/2] <= _S23i16[0];
			s23[mod*i+17] <= _S23i17[1];
			s23[mod*i+17+mod/2] <= _S23i17[0];
			s23[mod*i+18] <= _S23i18[1];
			s23[mod*i+18+mod/2] <= _S23i18[0];
			s23[mod*i+19] <= _S23i19[1];
			s23[mod*i+19+mod/2] <= _S23i19[0];
			s23[mod*i+20] <= _S23i20[1];
			s23[mod*i+20+mod/2] <= _S23i20[0];
			s23[mod*i+21] <= _S23i21[1];
			s23[mod*i+21+mod/2] <= _S23i21[0];
			s23[mod*i+22] <= _S23i22[1];
			s23[mod*i+22+mod/2] <= _S23i22[0];
			s23[mod*i+23] <= _S23i23[1];
			s23[mod*i+23+mod/2] <= _S23i23[0];
			s23[mod*i+24] <= _S23i24[1];
			s23[mod*i+24+mod/2] <= _S23i24[0];
			s23[mod*i+25] <= _S23i25[1];
			s23[mod*i+25+mod/2] <= _S23i25[0];
			s23[mod*i+26] <= _S23i26[1];
			s23[mod*i+26+mod/2] <= _S23i26[0];
			s23[mod*i+27] <= _S23i27[1];
			s23[mod*i+27+mod/2] <= _S23i27[0];
			s23[mod*i+28] <= _S23i28[1];
			s23[mod*i+28+mod/2] <= _S23i28[0];
			s23[mod*i+29] <= _S23i29[1];
			s23[mod*i+29+mod/2] <= _S23i29[0];
			s23[mod*i+30] <= _S23i30[1];
			s23[mod*i+30+mod/2] <= _S23i30[0];
			s23[mod*i+31] <= _S23i31[1];
			s23[mod*i+31+mod/2] <= _S23i31[0];
		end
	end
	p23.enq(1);
endrule
rule _Q65;
	p23.deq;
	let mod = 32;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S24i0 = min_max(pack(s23[mod*i+0]) , pack(s23[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S24i1 = min_max(pack(s23[mod*i+1]) , pack(s23[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S24i2 = min_max(pack(s23[mod*i+2]) , pack(s23[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S24i3 = min_max(pack(s23[mod*i+3]) , pack(s23[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S24i4 = min_max(pack(s23[mod*i+4]) , pack(s23[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S24i5 = min_max(pack(s23[mod*i+5]) , pack(s23[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S24i6 = min_max(pack(s23[mod*i+6]) , pack(s23[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S24i7 = min_max(pack(s23[mod*i+7]) , pack(s23[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S24i8 = min_max(pack(s23[mod*i+8]) , pack(s23[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S24i9 = min_max(pack(s23[mod*i+9]) , pack(s23[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S24i10 = min_max(pack(s23[mod*i+10]) , pack(s23[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S24i11 = min_max(pack(s23[mod*i+11]) , pack(s23[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S24i12 = min_max(pack(s23[mod*i+12]) , pack(s23[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S24i13 = min_max(pack(s23[mod*i+13]) , pack(s23[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S24i14 = min_max(pack(s23[mod*i+14]) , pack(s23[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S24i15 = min_max(pack(s23[mod*i+15]) , pack(s23[mod*i+15+mod/2]));
		if ((i/4)%2 == 0) begin
			s24[mod*i+0] <= _S24i0[0];
			s24[mod*i+0+mod/2] <= _S24i0[1];
			s24[mod*i+1] <= _S24i1[0];
			s24[mod*i+1+mod/2] <= _S24i1[1];
			s24[mod*i+2] <= _S24i2[0];
			s24[mod*i+2+mod/2] <= _S24i2[1];
			s24[mod*i+3] <= _S24i3[0];
			s24[mod*i+3+mod/2] <= _S24i3[1];
			s24[mod*i+4] <= _S24i4[0];
			s24[mod*i+4+mod/2] <= _S24i4[1];
			s24[mod*i+5] <= _S24i5[0];
			s24[mod*i+5+mod/2] <= _S24i5[1];
			s24[mod*i+6] <= _S24i6[0];
			s24[mod*i+6+mod/2] <= _S24i6[1];
			s24[mod*i+7] <= _S24i7[0];
			s24[mod*i+7+mod/2] <= _S24i7[1];
			s24[mod*i+8] <= _S24i8[0];
			s24[mod*i+8+mod/2] <= _S24i8[1];
			s24[mod*i+9] <= _S24i9[0];
			s24[mod*i+9+mod/2] <= _S24i9[1];
			s24[mod*i+10] <= _S24i10[0];
			s24[mod*i+10+mod/2] <= _S24i10[1];
			s24[mod*i+11] <= _S24i11[0];
			s24[mod*i+11+mod/2] <= _S24i11[1];
			s24[mod*i+12] <= _S24i12[0];
			s24[mod*i+12+mod/2] <= _S24i12[1];
			s24[mod*i+13] <= _S24i13[0];
			s24[mod*i+13+mod/2] <= _S24i13[1];
			s24[mod*i+14] <= _S24i14[0];
			s24[mod*i+14+mod/2] <= _S24i14[1];
			s24[mod*i+15] <= _S24i15[0];
			s24[mod*i+15+mod/2] <= _S24i15[1];
		end
		else begin
			s24[mod*i+0] <= _S24i0[1];
			s24[mod*i+0+mod/2] <= _S24i0[0];
			s24[mod*i+1] <= _S24i1[1];
			s24[mod*i+1+mod/2] <= _S24i1[0];
			s24[mod*i+2] <= _S24i2[1];
			s24[mod*i+2+mod/2] <= _S24i2[0];
			s24[mod*i+3] <= _S24i3[1];
			s24[mod*i+3+mod/2] <= _S24i3[0];
			s24[mod*i+4] <= _S24i4[1];
			s24[mod*i+4+mod/2] <= _S24i4[0];
			s24[mod*i+5] <= _S24i5[1];
			s24[mod*i+5+mod/2] <= _S24i5[0];
			s24[mod*i+6] <= _S24i6[1];
			s24[mod*i+6+mod/2] <= _S24i6[0];
			s24[mod*i+7] <= _S24i7[1];
			s24[mod*i+7+mod/2] <= _S24i7[0];
			s24[mod*i+8] <= _S24i8[1];
			s24[mod*i+8+mod/2] <= _S24i8[0];
			s24[mod*i+9] <= _S24i9[1];
			s24[mod*i+9+mod/2] <= _S24i9[0];
			s24[mod*i+10] <= _S24i10[1];
			s24[mod*i+10+mod/2] <= _S24i10[0];
			s24[mod*i+11] <= _S24i11[1];
			s24[mod*i+11+mod/2] <= _S24i11[0];
			s24[mod*i+12] <= _S24i12[1];
			s24[mod*i+12+mod/2] <= _S24i12[0];
			s24[mod*i+13] <= _S24i13[1];
			s24[mod*i+13+mod/2] <= _S24i13[0];
			s24[mod*i+14] <= _S24i14[1];
			s24[mod*i+14+mod/2] <= _S24i14[0];
			s24[mod*i+15] <= _S24i15[1];
			s24[mod*i+15+mod/2] <= _S24i15[0];
		end
	end
	p24.enq(1);
endrule
rule _Q64;
	p24.deq;
	let mod = 16;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S25i0 = min_max(pack(s24[mod*i+0]) , pack(s24[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S25i1 = min_max(pack(s24[mod*i+1]) , pack(s24[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S25i2 = min_max(pack(s24[mod*i+2]) , pack(s24[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S25i3 = min_max(pack(s24[mod*i+3]) , pack(s24[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S25i4 = min_max(pack(s24[mod*i+4]) , pack(s24[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S25i5 = min_max(pack(s24[mod*i+5]) , pack(s24[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S25i6 = min_max(pack(s24[mod*i+6]) , pack(s24[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S25i7 = min_max(pack(s24[mod*i+7]) , pack(s24[mod*i+7+mod/2]));
		if ((i/8)%2 == 0) begin
			s25[mod*i+0] <= _S25i0[0];
			s25[mod*i+0+mod/2] <= _S25i0[1];
			s25[mod*i+1] <= _S25i1[0];
			s25[mod*i+1+mod/2] <= _S25i1[1];
			s25[mod*i+2] <= _S25i2[0];
			s25[mod*i+2+mod/2] <= _S25i2[1];
			s25[mod*i+3] <= _S25i3[0];
			s25[mod*i+3+mod/2] <= _S25i3[1];
			s25[mod*i+4] <= _S25i4[0];
			s25[mod*i+4+mod/2] <= _S25i4[1];
			s25[mod*i+5] <= _S25i5[0];
			s25[mod*i+5+mod/2] <= _S25i5[1];
			s25[mod*i+6] <= _S25i6[0];
			s25[mod*i+6+mod/2] <= _S25i6[1];
			s25[mod*i+7] <= _S25i7[0];
			s25[mod*i+7+mod/2] <= _S25i7[1];
		end
		else begin
			s25[mod*i+0] <= _S25i0[1];
			s25[mod*i+0+mod/2] <= _S25i0[0];
			s25[mod*i+1] <= _S25i1[1];
			s25[mod*i+1+mod/2] <= _S25i1[0];
			s25[mod*i+2] <= _S25i2[1];
			s25[mod*i+2+mod/2] <= _S25i2[0];
			s25[mod*i+3] <= _S25i3[1];
			s25[mod*i+3+mod/2] <= _S25i3[0];
			s25[mod*i+4] <= _S25i4[1];
			s25[mod*i+4+mod/2] <= _S25i4[0];
			s25[mod*i+5] <= _S25i5[1];
			s25[mod*i+5+mod/2] <= _S25i5[0];
			s25[mod*i+6] <= _S25i6[1];
			s25[mod*i+6+mod/2] <= _S25i6[0];
			s25[mod*i+7] <= _S25i7[1];
			s25[mod*i+7+mod/2] <= _S25i7[0];
		end
	end
	p25.enq(1);
endrule
rule _Q63;
	p25.deq;
	let mod = 8;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S26i0 = min_max(pack(s25[mod*i+0]) , pack(s25[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S26i1 = min_max(pack(s25[mod*i+1]) , pack(s25[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S26i2 = min_max(pack(s25[mod*i+2]) , pack(s25[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S26i3 = min_max(pack(s25[mod*i+3]) , pack(s25[mod*i+3+mod/2]));
		if ((i/16)%2 == 0) begin
			s26[mod*i+0] <= _S26i0[0];
			s26[mod*i+0+mod/2] <= _S26i0[1];
			s26[mod*i+1] <= _S26i1[0];
			s26[mod*i+1+mod/2] <= _S26i1[1];
			s26[mod*i+2] <= _S26i2[0];
			s26[mod*i+2+mod/2] <= _S26i2[1];
			s26[mod*i+3] <= _S26i3[0];
			s26[mod*i+3+mod/2] <= _S26i3[1];
		end
		else begin
			s26[mod*i+0] <= _S26i0[1];
			s26[mod*i+0+mod/2] <= _S26i0[0];
			s26[mod*i+1] <= _S26i1[1];
			s26[mod*i+1+mod/2] <= _S26i1[0];
			s26[mod*i+2] <= _S26i2[1];
			s26[mod*i+2+mod/2] <= _S26i2[0];
			s26[mod*i+3] <= _S26i3[1];
			s26[mod*i+3+mod/2] <= _S26i3[0];
		end
	end
	p26.enq(1);
endrule
rule _Q62;
	p26.deq;
	let mod = 4;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S27i0 = min_max(pack(s26[mod*i+0]) , pack(s26[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S27i1 = min_max(pack(s26[mod*i+1]) , pack(s26[mod*i+1+mod/2]));
		if ((i/32)%2 == 0) begin
			s27[mod*i+0] <= _S27i0[0];
			s27[mod*i+0+mod/2] <= _S27i0[1];
			s27[mod*i+1] <= _S27i1[0];
			s27[mod*i+1+mod/2] <= _S27i1[1];
		end
		else begin
			s27[mod*i+0] <= _S27i0[1];
			s27[mod*i+0+mod/2] <= _S27i0[0];
			s27[mod*i+1] <= _S27i1[1];
			s27[mod*i+1+mod/2] <= _S27i1[0];
		end
	end
	p27.enq(1);
endrule
rule _Q61;
	p27.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S28i0 = min_max(pack(s27[mod*i+0]) , pack(s27[mod*i+0+mod/2]));
		if ((i/64)%2 == 0) begin
			s28[mod*i+0] <= _S28i0[0];
			s28[mod*i+0+mod/2] <= _S28i0[1];
		end
		else begin
			s28[mod*i+0] <= _S28i0[1];
			s28[mod*i+0+mod/2] <= _S28i0[0];
		end
	end
	p28.enq(1);
endrule
rule _Q78;
	p28.deq;
	let mod = 256;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S29i0 = min_max(pack(s28[mod*i+0]) , pack(s28[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S29i1 = min_max(pack(s28[mod*i+1]) , pack(s28[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S29i2 = min_max(pack(s28[mod*i+2]) , pack(s28[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S29i3 = min_max(pack(s28[mod*i+3]) , pack(s28[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S29i4 = min_max(pack(s28[mod*i+4]) , pack(s28[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S29i5 = min_max(pack(s28[mod*i+5]) , pack(s28[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S29i6 = min_max(pack(s28[mod*i+6]) , pack(s28[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S29i7 = min_max(pack(s28[mod*i+7]) , pack(s28[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S29i8 = min_max(pack(s28[mod*i+8]) , pack(s28[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S29i9 = min_max(pack(s28[mod*i+9]) , pack(s28[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S29i10 = min_max(pack(s28[mod*i+10]) , pack(s28[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S29i11 = min_max(pack(s28[mod*i+11]) , pack(s28[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S29i12 = min_max(pack(s28[mod*i+12]) , pack(s28[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S29i13 = min_max(pack(s28[mod*i+13]) , pack(s28[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S29i14 = min_max(pack(s28[mod*i+14]) , pack(s28[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S29i15 = min_max(pack(s28[mod*i+15]) , pack(s28[mod*i+15+mod/2]));
			 Vector#(2, Int#(32)) _S29i16 = min_max(pack(s28[mod*i+16]) , pack(s28[mod*i+16+mod/2]));
			 Vector#(2, Int#(32)) _S29i17 = min_max(pack(s28[mod*i+17]) , pack(s28[mod*i+17+mod/2]));
			 Vector#(2, Int#(32)) _S29i18 = min_max(pack(s28[mod*i+18]) , pack(s28[mod*i+18+mod/2]));
			 Vector#(2, Int#(32)) _S29i19 = min_max(pack(s28[mod*i+19]) , pack(s28[mod*i+19+mod/2]));
			 Vector#(2, Int#(32)) _S29i20 = min_max(pack(s28[mod*i+20]) , pack(s28[mod*i+20+mod/2]));
			 Vector#(2, Int#(32)) _S29i21 = min_max(pack(s28[mod*i+21]) , pack(s28[mod*i+21+mod/2]));
			 Vector#(2, Int#(32)) _S29i22 = min_max(pack(s28[mod*i+22]) , pack(s28[mod*i+22+mod/2]));
			 Vector#(2, Int#(32)) _S29i23 = min_max(pack(s28[mod*i+23]) , pack(s28[mod*i+23+mod/2]));
			 Vector#(2, Int#(32)) _S29i24 = min_max(pack(s28[mod*i+24]) , pack(s28[mod*i+24+mod/2]));
			 Vector#(2, Int#(32)) _S29i25 = min_max(pack(s28[mod*i+25]) , pack(s28[mod*i+25+mod/2]));
			 Vector#(2, Int#(32)) _S29i26 = min_max(pack(s28[mod*i+26]) , pack(s28[mod*i+26+mod/2]));
			 Vector#(2, Int#(32)) _S29i27 = min_max(pack(s28[mod*i+27]) , pack(s28[mod*i+27+mod/2]));
			 Vector#(2, Int#(32)) _S29i28 = min_max(pack(s28[mod*i+28]) , pack(s28[mod*i+28+mod/2]));
			 Vector#(2, Int#(32)) _S29i29 = min_max(pack(s28[mod*i+29]) , pack(s28[mod*i+29+mod/2]));
			 Vector#(2, Int#(32)) _S29i30 = min_max(pack(s28[mod*i+30]) , pack(s28[mod*i+30+mod/2]));
			 Vector#(2, Int#(32)) _S29i31 = min_max(pack(s28[mod*i+31]) , pack(s28[mod*i+31+mod/2]));
			 Vector#(2, Int#(32)) _S29i32 = min_max(pack(s28[mod*i+32]) , pack(s28[mod*i+32+mod/2]));
			 Vector#(2, Int#(32)) _S29i33 = min_max(pack(s28[mod*i+33]) , pack(s28[mod*i+33+mod/2]));
			 Vector#(2, Int#(32)) _S29i34 = min_max(pack(s28[mod*i+34]) , pack(s28[mod*i+34+mod/2]));
			 Vector#(2, Int#(32)) _S29i35 = min_max(pack(s28[mod*i+35]) , pack(s28[mod*i+35+mod/2]));
			 Vector#(2, Int#(32)) _S29i36 = min_max(pack(s28[mod*i+36]) , pack(s28[mod*i+36+mod/2]));
			 Vector#(2, Int#(32)) _S29i37 = min_max(pack(s28[mod*i+37]) , pack(s28[mod*i+37+mod/2]));
			 Vector#(2, Int#(32)) _S29i38 = min_max(pack(s28[mod*i+38]) , pack(s28[mod*i+38+mod/2]));
			 Vector#(2, Int#(32)) _S29i39 = min_max(pack(s28[mod*i+39]) , pack(s28[mod*i+39+mod/2]));
			 Vector#(2, Int#(32)) _S29i40 = min_max(pack(s28[mod*i+40]) , pack(s28[mod*i+40+mod/2]));
			 Vector#(2, Int#(32)) _S29i41 = min_max(pack(s28[mod*i+41]) , pack(s28[mod*i+41+mod/2]));
			 Vector#(2, Int#(32)) _S29i42 = min_max(pack(s28[mod*i+42]) , pack(s28[mod*i+42+mod/2]));
			 Vector#(2, Int#(32)) _S29i43 = min_max(pack(s28[mod*i+43]) , pack(s28[mod*i+43+mod/2]));
			 Vector#(2, Int#(32)) _S29i44 = min_max(pack(s28[mod*i+44]) , pack(s28[mod*i+44+mod/2]));
			 Vector#(2, Int#(32)) _S29i45 = min_max(pack(s28[mod*i+45]) , pack(s28[mod*i+45+mod/2]));
			 Vector#(2, Int#(32)) _S29i46 = min_max(pack(s28[mod*i+46]) , pack(s28[mod*i+46+mod/2]));
			 Vector#(2, Int#(32)) _S29i47 = min_max(pack(s28[mod*i+47]) , pack(s28[mod*i+47+mod/2]));
			 Vector#(2, Int#(32)) _S29i48 = min_max(pack(s28[mod*i+48]) , pack(s28[mod*i+48+mod/2]));
			 Vector#(2, Int#(32)) _S29i49 = min_max(pack(s28[mod*i+49]) , pack(s28[mod*i+49+mod/2]));
			 Vector#(2, Int#(32)) _S29i50 = min_max(pack(s28[mod*i+50]) , pack(s28[mod*i+50+mod/2]));
			 Vector#(2, Int#(32)) _S29i51 = min_max(pack(s28[mod*i+51]) , pack(s28[mod*i+51+mod/2]));
			 Vector#(2, Int#(32)) _S29i52 = min_max(pack(s28[mod*i+52]) , pack(s28[mod*i+52+mod/2]));
			 Vector#(2, Int#(32)) _S29i53 = min_max(pack(s28[mod*i+53]) , pack(s28[mod*i+53+mod/2]));
			 Vector#(2, Int#(32)) _S29i54 = min_max(pack(s28[mod*i+54]) , pack(s28[mod*i+54+mod/2]));
			 Vector#(2, Int#(32)) _S29i55 = min_max(pack(s28[mod*i+55]) , pack(s28[mod*i+55+mod/2]));
			 Vector#(2, Int#(32)) _S29i56 = min_max(pack(s28[mod*i+56]) , pack(s28[mod*i+56+mod/2]));
			 Vector#(2, Int#(32)) _S29i57 = min_max(pack(s28[mod*i+57]) , pack(s28[mod*i+57+mod/2]));
			 Vector#(2, Int#(32)) _S29i58 = min_max(pack(s28[mod*i+58]) , pack(s28[mod*i+58+mod/2]));
			 Vector#(2, Int#(32)) _S29i59 = min_max(pack(s28[mod*i+59]) , pack(s28[mod*i+59+mod/2]));
			 Vector#(2, Int#(32)) _S29i60 = min_max(pack(s28[mod*i+60]) , pack(s28[mod*i+60+mod/2]));
			 Vector#(2, Int#(32)) _S29i61 = min_max(pack(s28[mod*i+61]) , pack(s28[mod*i+61+mod/2]));
			 Vector#(2, Int#(32)) _S29i62 = min_max(pack(s28[mod*i+62]) , pack(s28[mod*i+62+mod/2]));
			 Vector#(2, Int#(32)) _S29i63 = min_max(pack(s28[mod*i+63]) , pack(s28[mod*i+63+mod/2]));
			 Vector#(2, Int#(32)) _S29i64 = min_max(pack(s28[mod*i+64]) , pack(s28[mod*i+64+mod/2]));
			 Vector#(2, Int#(32)) _S29i65 = min_max(pack(s28[mod*i+65]) , pack(s28[mod*i+65+mod/2]));
			 Vector#(2, Int#(32)) _S29i66 = min_max(pack(s28[mod*i+66]) , pack(s28[mod*i+66+mod/2]));
			 Vector#(2, Int#(32)) _S29i67 = min_max(pack(s28[mod*i+67]) , pack(s28[mod*i+67+mod/2]));
			 Vector#(2, Int#(32)) _S29i68 = min_max(pack(s28[mod*i+68]) , pack(s28[mod*i+68+mod/2]));
			 Vector#(2, Int#(32)) _S29i69 = min_max(pack(s28[mod*i+69]) , pack(s28[mod*i+69+mod/2]));
			 Vector#(2, Int#(32)) _S29i70 = min_max(pack(s28[mod*i+70]) , pack(s28[mod*i+70+mod/2]));
			 Vector#(2, Int#(32)) _S29i71 = min_max(pack(s28[mod*i+71]) , pack(s28[mod*i+71+mod/2]));
			 Vector#(2, Int#(32)) _S29i72 = min_max(pack(s28[mod*i+72]) , pack(s28[mod*i+72+mod/2]));
			 Vector#(2, Int#(32)) _S29i73 = min_max(pack(s28[mod*i+73]) , pack(s28[mod*i+73+mod/2]));
			 Vector#(2, Int#(32)) _S29i74 = min_max(pack(s28[mod*i+74]) , pack(s28[mod*i+74+mod/2]));
			 Vector#(2, Int#(32)) _S29i75 = min_max(pack(s28[mod*i+75]) , pack(s28[mod*i+75+mod/2]));
			 Vector#(2, Int#(32)) _S29i76 = min_max(pack(s28[mod*i+76]) , pack(s28[mod*i+76+mod/2]));
			 Vector#(2, Int#(32)) _S29i77 = min_max(pack(s28[mod*i+77]) , pack(s28[mod*i+77+mod/2]));
			 Vector#(2, Int#(32)) _S29i78 = min_max(pack(s28[mod*i+78]) , pack(s28[mod*i+78+mod/2]));
			 Vector#(2, Int#(32)) _S29i79 = min_max(pack(s28[mod*i+79]) , pack(s28[mod*i+79+mod/2]));
			 Vector#(2, Int#(32)) _S29i80 = min_max(pack(s28[mod*i+80]) , pack(s28[mod*i+80+mod/2]));
			 Vector#(2, Int#(32)) _S29i81 = min_max(pack(s28[mod*i+81]) , pack(s28[mod*i+81+mod/2]));
			 Vector#(2, Int#(32)) _S29i82 = min_max(pack(s28[mod*i+82]) , pack(s28[mod*i+82+mod/2]));
			 Vector#(2, Int#(32)) _S29i83 = min_max(pack(s28[mod*i+83]) , pack(s28[mod*i+83+mod/2]));
			 Vector#(2, Int#(32)) _S29i84 = min_max(pack(s28[mod*i+84]) , pack(s28[mod*i+84+mod/2]));
			 Vector#(2, Int#(32)) _S29i85 = min_max(pack(s28[mod*i+85]) , pack(s28[mod*i+85+mod/2]));
			 Vector#(2, Int#(32)) _S29i86 = min_max(pack(s28[mod*i+86]) , pack(s28[mod*i+86+mod/2]));
			 Vector#(2, Int#(32)) _S29i87 = min_max(pack(s28[mod*i+87]) , pack(s28[mod*i+87+mod/2]));
			 Vector#(2, Int#(32)) _S29i88 = min_max(pack(s28[mod*i+88]) , pack(s28[mod*i+88+mod/2]));
			 Vector#(2, Int#(32)) _S29i89 = min_max(pack(s28[mod*i+89]) , pack(s28[mod*i+89+mod/2]));
			 Vector#(2, Int#(32)) _S29i90 = min_max(pack(s28[mod*i+90]) , pack(s28[mod*i+90+mod/2]));
			 Vector#(2, Int#(32)) _S29i91 = min_max(pack(s28[mod*i+91]) , pack(s28[mod*i+91+mod/2]));
			 Vector#(2, Int#(32)) _S29i92 = min_max(pack(s28[mod*i+92]) , pack(s28[mod*i+92+mod/2]));
			 Vector#(2, Int#(32)) _S29i93 = min_max(pack(s28[mod*i+93]) , pack(s28[mod*i+93+mod/2]));
			 Vector#(2, Int#(32)) _S29i94 = min_max(pack(s28[mod*i+94]) , pack(s28[mod*i+94+mod/2]));
			 Vector#(2, Int#(32)) _S29i95 = min_max(pack(s28[mod*i+95]) , pack(s28[mod*i+95+mod/2]));
			 Vector#(2, Int#(32)) _S29i96 = min_max(pack(s28[mod*i+96]) , pack(s28[mod*i+96+mod/2]));
			 Vector#(2, Int#(32)) _S29i97 = min_max(pack(s28[mod*i+97]) , pack(s28[mod*i+97+mod/2]));
			 Vector#(2, Int#(32)) _S29i98 = min_max(pack(s28[mod*i+98]) , pack(s28[mod*i+98+mod/2]));
			 Vector#(2, Int#(32)) _S29i99 = min_max(pack(s28[mod*i+99]) , pack(s28[mod*i+99+mod/2]));
			 Vector#(2, Int#(32)) _S29i100 = min_max(pack(s28[mod*i+100]) , pack(s28[mod*i+100+mod/2]));
			 Vector#(2, Int#(32)) _S29i101 = min_max(pack(s28[mod*i+101]) , pack(s28[mod*i+101+mod/2]));
			 Vector#(2, Int#(32)) _S29i102 = min_max(pack(s28[mod*i+102]) , pack(s28[mod*i+102+mod/2]));
			 Vector#(2, Int#(32)) _S29i103 = min_max(pack(s28[mod*i+103]) , pack(s28[mod*i+103+mod/2]));
			 Vector#(2, Int#(32)) _S29i104 = min_max(pack(s28[mod*i+104]) , pack(s28[mod*i+104+mod/2]));
			 Vector#(2, Int#(32)) _S29i105 = min_max(pack(s28[mod*i+105]) , pack(s28[mod*i+105+mod/2]));
			 Vector#(2, Int#(32)) _S29i106 = min_max(pack(s28[mod*i+106]) , pack(s28[mod*i+106+mod/2]));
			 Vector#(2, Int#(32)) _S29i107 = min_max(pack(s28[mod*i+107]) , pack(s28[mod*i+107+mod/2]));
			 Vector#(2, Int#(32)) _S29i108 = min_max(pack(s28[mod*i+108]) , pack(s28[mod*i+108+mod/2]));
			 Vector#(2, Int#(32)) _S29i109 = min_max(pack(s28[mod*i+109]) , pack(s28[mod*i+109+mod/2]));
			 Vector#(2, Int#(32)) _S29i110 = min_max(pack(s28[mod*i+110]) , pack(s28[mod*i+110+mod/2]));
			 Vector#(2, Int#(32)) _S29i111 = min_max(pack(s28[mod*i+111]) , pack(s28[mod*i+111+mod/2]));
			 Vector#(2, Int#(32)) _S29i112 = min_max(pack(s28[mod*i+112]) , pack(s28[mod*i+112+mod/2]));
			 Vector#(2, Int#(32)) _S29i113 = min_max(pack(s28[mod*i+113]) , pack(s28[mod*i+113+mod/2]));
			 Vector#(2, Int#(32)) _S29i114 = min_max(pack(s28[mod*i+114]) , pack(s28[mod*i+114+mod/2]));
			 Vector#(2, Int#(32)) _S29i115 = min_max(pack(s28[mod*i+115]) , pack(s28[mod*i+115+mod/2]));
			 Vector#(2, Int#(32)) _S29i116 = min_max(pack(s28[mod*i+116]) , pack(s28[mod*i+116+mod/2]));
			 Vector#(2, Int#(32)) _S29i117 = min_max(pack(s28[mod*i+117]) , pack(s28[mod*i+117+mod/2]));
			 Vector#(2, Int#(32)) _S29i118 = min_max(pack(s28[mod*i+118]) , pack(s28[mod*i+118+mod/2]));
			 Vector#(2, Int#(32)) _S29i119 = min_max(pack(s28[mod*i+119]) , pack(s28[mod*i+119+mod/2]));
			 Vector#(2, Int#(32)) _S29i120 = min_max(pack(s28[mod*i+120]) , pack(s28[mod*i+120+mod/2]));
			 Vector#(2, Int#(32)) _S29i121 = min_max(pack(s28[mod*i+121]) , pack(s28[mod*i+121+mod/2]));
			 Vector#(2, Int#(32)) _S29i122 = min_max(pack(s28[mod*i+122]) , pack(s28[mod*i+122+mod/2]));
			 Vector#(2, Int#(32)) _S29i123 = min_max(pack(s28[mod*i+123]) , pack(s28[mod*i+123+mod/2]));
			 Vector#(2, Int#(32)) _S29i124 = min_max(pack(s28[mod*i+124]) , pack(s28[mod*i+124+mod/2]));
			 Vector#(2, Int#(32)) _S29i125 = min_max(pack(s28[mod*i+125]) , pack(s28[mod*i+125+mod/2]));
			 Vector#(2, Int#(32)) _S29i126 = min_max(pack(s28[mod*i+126]) , pack(s28[mod*i+126+mod/2]));
			 Vector#(2, Int#(32)) _S29i127 = min_max(pack(s28[mod*i+127]) , pack(s28[mod*i+127+mod/2]));
		if ((i/1)%2 == 0) begin
			s29[mod*i+0] <= _S29i0[0];
			s29[mod*i+0+mod/2] <= _S29i0[1];
			s29[mod*i+1] <= _S29i1[0];
			s29[mod*i+1+mod/2] <= _S29i1[1];
			s29[mod*i+2] <= _S29i2[0];
			s29[mod*i+2+mod/2] <= _S29i2[1];
			s29[mod*i+3] <= _S29i3[0];
			s29[mod*i+3+mod/2] <= _S29i3[1];
			s29[mod*i+4] <= _S29i4[0];
			s29[mod*i+4+mod/2] <= _S29i4[1];
			s29[mod*i+5] <= _S29i5[0];
			s29[mod*i+5+mod/2] <= _S29i5[1];
			s29[mod*i+6] <= _S29i6[0];
			s29[mod*i+6+mod/2] <= _S29i6[1];
			s29[mod*i+7] <= _S29i7[0];
			s29[mod*i+7+mod/2] <= _S29i7[1];
			s29[mod*i+8] <= _S29i8[0];
			s29[mod*i+8+mod/2] <= _S29i8[1];
			s29[mod*i+9] <= _S29i9[0];
			s29[mod*i+9+mod/2] <= _S29i9[1];
			s29[mod*i+10] <= _S29i10[0];
			s29[mod*i+10+mod/2] <= _S29i10[1];
			s29[mod*i+11] <= _S29i11[0];
			s29[mod*i+11+mod/2] <= _S29i11[1];
			s29[mod*i+12] <= _S29i12[0];
			s29[mod*i+12+mod/2] <= _S29i12[1];
			s29[mod*i+13] <= _S29i13[0];
			s29[mod*i+13+mod/2] <= _S29i13[1];
			s29[mod*i+14] <= _S29i14[0];
			s29[mod*i+14+mod/2] <= _S29i14[1];
			s29[mod*i+15] <= _S29i15[0];
			s29[mod*i+15+mod/2] <= _S29i15[1];
			s29[mod*i+16] <= _S29i16[0];
			s29[mod*i+16+mod/2] <= _S29i16[1];
			s29[mod*i+17] <= _S29i17[0];
			s29[mod*i+17+mod/2] <= _S29i17[1];
			s29[mod*i+18] <= _S29i18[0];
			s29[mod*i+18+mod/2] <= _S29i18[1];
			s29[mod*i+19] <= _S29i19[0];
			s29[mod*i+19+mod/2] <= _S29i19[1];
			s29[mod*i+20] <= _S29i20[0];
			s29[mod*i+20+mod/2] <= _S29i20[1];
			s29[mod*i+21] <= _S29i21[0];
			s29[mod*i+21+mod/2] <= _S29i21[1];
			s29[mod*i+22] <= _S29i22[0];
			s29[mod*i+22+mod/2] <= _S29i22[1];
			s29[mod*i+23] <= _S29i23[0];
			s29[mod*i+23+mod/2] <= _S29i23[1];
			s29[mod*i+24] <= _S29i24[0];
			s29[mod*i+24+mod/2] <= _S29i24[1];
			s29[mod*i+25] <= _S29i25[0];
			s29[mod*i+25+mod/2] <= _S29i25[1];
			s29[mod*i+26] <= _S29i26[0];
			s29[mod*i+26+mod/2] <= _S29i26[1];
			s29[mod*i+27] <= _S29i27[0];
			s29[mod*i+27+mod/2] <= _S29i27[1];
			s29[mod*i+28] <= _S29i28[0];
			s29[mod*i+28+mod/2] <= _S29i28[1];
			s29[mod*i+29] <= _S29i29[0];
			s29[mod*i+29+mod/2] <= _S29i29[1];
			s29[mod*i+30] <= _S29i30[0];
			s29[mod*i+30+mod/2] <= _S29i30[1];
			s29[mod*i+31] <= _S29i31[0];
			s29[mod*i+31+mod/2] <= _S29i31[1];
			s29[mod*i+32] <= _S29i32[0];
			s29[mod*i+32+mod/2] <= _S29i32[1];
			s29[mod*i+33] <= _S29i33[0];
			s29[mod*i+33+mod/2] <= _S29i33[1];
			s29[mod*i+34] <= _S29i34[0];
			s29[mod*i+34+mod/2] <= _S29i34[1];
			s29[mod*i+35] <= _S29i35[0];
			s29[mod*i+35+mod/2] <= _S29i35[1];
			s29[mod*i+36] <= _S29i36[0];
			s29[mod*i+36+mod/2] <= _S29i36[1];
			s29[mod*i+37] <= _S29i37[0];
			s29[mod*i+37+mod/2] <= _S29i37[1];
			s29[mod*i+38] <= _S29i38[0];
			s29[mod*i+38+mod/2] <= _S29i38[1];
			s29[mod*i+39] <= _S29i39[0];
			s29[mod*i+39+mod/2] <= _S29i39[1];
			s29[mod*i+40] <= _S29i40[0];
			s29[mod*i+40+mod/2] <= _S29i40[1];
			s29[mod*i+41] <= _S29i41[0];
			s29[mod*i+41+mod/2] <= _S29i41[1];
			s29[mod*i+42] <= _S29i42[0];
			s29[mod*i+42+mod/2] <= _S29i42[1];
			s29[mod*i+43] <= _S29i43[0];
			s29[mod*i+43+mod/2] <= _S29i43[1];
			s29[mod*i+44] <= _S29i44[0];
			s29[mod*i+44+mod/2] <= _S29i44[1];
			s29[mod*i+45] <= _S29i45[0];
			s29[mod*i+45+mod/2] <= _S29i45[1];
			s29[mod*i+46] <= _S29i46[0];
			s29[mod*i+46+mod/2] <= _S29i46[1];
			s29[mod*i+47] <= _S29i47[0];
			s29[mod*i+47+mod/2] <= _S29i47[1];
			s29[mod*i+48] <= _S29i48[0];
			s29[mod*i+48+mod/2] <= _S29i48[1];
			s29[mod*i+49] <= _S29i49[0];
			s29[mod*i+49+mod/2] <= _S29i49[1];
			s29[mod*i+50] <= _S29i50[0];
			s29[mod*i+50+mod/2] <= _S29i50[1];
			s29[mod*i+51] <= _S29i51[0];
			s29[mod*i+51+mod/2] <= _S29i51[1];
			s29[mod*i+52] <= _S29i52[0];
			s29[mod*i+52+mod/2] <= _S29i52[1];
			s29[mod*i+53] <= _S29i53[0];
			s29[mod*i+53+mod/2] <= _S29i53[1];
			s29[mod*i+54] <= _S29i54[0];
			s29[mod*i+54+mod/2] <= _S29i54[1];
			s29[mod*i+55] <= _S29i55[0];
			s29[mod*i+55+mod/2] <= _S29i55[1];
			s29[mod*i+56] <= _S29i56[0];
			s29[mod*i+56+mod/2] <= _S29i56[1];
			s29[mod*i+57] <= _S29i57[0];
			s29[mod*i+57+mod/2] <= _S29i57[1];
			s29[mod*i+58] <= _S29i58[0];
			s29[mod*i+58+mod/2] <= _S29i58[1];
			s29[mod*i+59] <= _S29i59[0];
			s29[mod*i+59+mod/2] <= _S29i59[1];
			s29[mod*i+60] <= _S29i60[0];
			s29[mod*i+60+mod/2] <= _S29i60[1];
			s29[mod*i+61] <= _S29i61[0];
			s29[mod*i+61+mod/2] <= _S29i61[1];
			s29[mod*i+62] <= _S29i62[0];
			s29[mod*i+62+mod/2] <= _S29i62[1];
			s29[mod*i+63] <= _S29i63[0];
			s29[mod*i+63+mod/2] <= _S29i63[1];
			s29[mod*i+64] <= _S29i64[0];
			s29[mod*i+64+mod/2] <= _S29i64[1];
			s29[mod*i+65] <= _S29i65[0];
			s29[mod*i+65+mod/2] <= _S29i65[1];
			s29[mod*i+66] <= _S29i66[0];
			s29[mod*i+66+mod/2] <= _S29i66[1];
			s29[mod*i+67] <= _S29i67[0];
			s29[mod*i+67+mod/2] <= _S29i67[1];
			s29[mod*i+68] <= _S29i68[0];
			s29[mod*i+68+mod/2] <= _S29i68[1];
			s29[mod*i+69] <= _S29i69[0];
			s29[mod*i+69+mod/2] <= _S29i69[1];
			s29[mod*i+70] <= _S29i70[0];
			s29[mod*i+70+mod/2] <= _S29i70[1];
			s29[mod*i+71] <= _S29i71[0];
			s29[mod*i+71+mod/2] <= _S29i71[1];
			s29[mod*i+72] <= _S29i72[0];
			s29[mod*i+72+mod/2] <= _S29i72[1];
			s29[mod*i+73] <= _S29i73[0];
			s29[mod*i+73+mod/2] <= _S29i73[1];
			s29[mod*i+74] <= _S29i74[0];
			s29[mod*i+74+mod/2] <= _S29i74[1];
			s29[mod*i+75] <= _S29i75[0];
			s29[mod*i+75+mod/2] <= _S29i75[1];
			s29[mod*i+76] <= _S29i76[0];
			s29[mod*i+76+mod/2] <= _S29i76[1];
			s29[mod*i+77] <= _S29i77[0];
			s29[mod*i+77+mod/2] <= _S29i77[1];
			s29[mod*i+78] <= _S29i78[0];
			s29[mod*i+78+mod/2] <= _S29i78[1];
			s29[mod*i+79] <= _S29i79[0];
			s29[mod*i+79+mod/2] <= _S29i79[1];
			s29[mod*i+80] <= _S29i80[0];
			s29[mod*i+80+mod/2] <= _S29i80[1];
			s29[mod*i+81] <= _S29i81[0];
			s29[mod*i+81+mod/2] <= _S29i81[1];
			s29[mod*i+82] <= _S29i82[0];
			s29[mod*i+82+mod/2] <= _S29i82[1];
			s29[mod*i+83] <= _S29i83[0];
			s29[mod*i+83+mod/2] <= _S29i83[1];
			s29[mod*i+84] <= _S29i84[0];
			s29[mod*i+84+mod/2] <= _S29i84[1];
			s29[mod*i+85] <= _S29i85[0];
			s29[mod*i+85+mod/2] <= _S29i85[1];
			s29[mod*i+86] <= _S29i86[0];
			s29[mod*i+86+mod/2] <= _S29i86[1];
			s29[mod*i+87] <= _S29i87[0];
			s29[mod*i+87+mod/2] <= _S29i87[1];
			s29[mod*i+88] <= _S29i88[0];
			s29[mod*i+88+mod/2] <= _S29i88[1];
			s29[mod*i+89] <= _S29i89[0];
			s29[mod*i+89+mod/2] <= _S29i89[1];
			s29[mod*i+90] <= _S29i90[0];
			s29[mod*i+90+mod/2] <= _S29i90[1];
			s29[mod*i+91] <= _S29i91[0];
			s29[mod*i+91+mod/2] <= _S29i91[1];
			s29[mod*i+92] <= _S29i92[0];
			s29[mod*i+92+mod/2] <= _S29i92[1];
			s29[mod*i+93] <= _S29i93[0];
			s29[mod*i+93+mod/2] <= _S29i93[1];
			s29[mod*i+94] <= _S29i94[0];
			s29[mod*i+94+mod/2] <= _S29i94[1];
			s29[mod*i+95] <= _S29i95[0];
			s29[mod*i+95+mod/2] <= _S29i95[1];
			s29[mod*i+96] <= _S29i96[0];
			s29[mod*i+96+mod/2] <= _S29i96[1];
			s29[mod*i+97] <= _S29i97[0];
			s29[mod*i+97+mod/2] <= _S29i97[1];
			s29[mod*i+98] <= _S29i98[0];
			s29[mod*i+98+mod/2] <= _S29i98[1];
			s29[mod*i+99] <= _S29i99[0];
			s29[mod*i+99+mod/2] <= _S29i99[1];
			s29[mod*i+100] <= _S29i100[0];
			s29[mod*i+100+mod/2] <= _S29i100[1];
			s29[mod*i+101] <= _S29i101[0];
			s29[mod*i+101+mod/2] <= _S29i101[1];
			s29[mod*i+102] <= _S29i102[0];
			s29[mod*i+102+mod/2] <= _S29i102[1];
			s29[mod*i+103] <= _S29i103[0];
			s29[mod*i+103+mod/2] <= _S29i103[1];
			s29[mod*i+104] <= _S29i104[0];
			s29[mod*i+104+mod/2] <= _S29i104[1];
			s29[mod*i+105] <= _S29i105[0];
			s29[mod*i+105+mod/2] <= _S29i105[1];
			s29[mod*i+106] <= _S29i106[0];
			s29[mod*i+106+mod/2] <= _S29i106[1];
			s29[mod*i+107] <= _S29i107[0];
			s29[mod*i+107+mod/2] <= _S29i107[1];
			s29[mod*i+108] <= _S29i108[0];
			s29[mod*i+108+mod/2] <= _S29i108[1];
			s29[mod*i+109] <= _S29i109[0];
			s29[mod*i+109+mod/2] <= _S29i109[1];
			s29[mod*i+110] <= _S29i110[0];
			s29[mod*i+110+mod/2] <= _S29i110[1];
			s29[mod*i+111] <= _S29i111[0];
			s29[mod*i+111+mod/2] <= _S29i111[1];
			s29[mod*i+112] <= _S29i112[0];
			s29[mod*i+112+mod/2] <= _S29i112[1];
			s29[mod*i+113] <= _S29i113[0];
			s29[mod*i+113+mod/2] <= _S29i113[1];
			s29[mod*i+114] <= _S29i114[0];
			s29[mod*i+114+mod/2] <= _S29i114[1];
			s29[mod*i+115] <= _S29i115[0];
			s29[mod*i+115+mod/2] <= _S29i115[1];
			s29[mod*i+116] <= _S29i116[0];
			s29[mod*i+116+mod/2] <= _S29i116[1];
			s29[mod*i+117] <= _S29i117[0];
			s29[mod*i+117+mod/2] <= _S29i117[1];
			s29[mod*i+118] <= _S29i118[0];
			s29[mod*i+118+mod/2] <= _S29i118[1];
			s29[mod*i+119] <= _S29i119[0];
			s29[mod*i+119+mod/2] <= _S29i119[1];
			s29[mod*i+120] <= _S29i120[0];
			s29[mod*i+120+mod/2] <= _S29i120[1];
			s29[mod*i+121] <= _S29i121[0];
			s29[mod*i+121+mod/2] <= _S29i121[1];
			s29[mod*i+122] <= _S29i122[0];
			s29[mod*i+122+mod/2] <= _S29i122[1];
			s29[mod*i+123] <= _S29i123[0];
			s29[mod*i+123+mod/2] <= _S29i123[1];
			s29[mod*i+124] <= _S29i124[0];
			s29[mod*i+124+mod/2] <= _S29i124[1];
			s29[mod*i+125] <= _S29i125[0];
			s29[mod*i+125+mod/2] <= _S29i125[1];
			s29[mod*i+126] <= _S29i126[0];
			s29[mod*i+126+mod/2] <= _S29i126[1];
			s29[mod*i+127] <= _S29i127[0];
			s29[mod*i+127+mod/2] <= _S29i127[1];
		end
		else begin
			s29[mod*i+0] <= _S29i0[1];
			s29[mod*i+0+mod/2] <= _S29i0[0];
			s29[mod*i+1] <= _S29i1[1];
			s29[mod*i+1+mod/2] <= _S29i1[0];
			s29[mod*i+2] <= _S29i2[1];
			s29[mod*i+2+mod/2] <= _S29i2[0];
			s29[mod*i+3] <= _S29i3[1];
			s29[mod*i+3+mod/2] <= _S29i3[0];
			s29[mod*i+4] <= _S29i4[1];
			s29[mod*i+4+mod/2] <= _S29i4[0];
			s29[mod*i+5] <= _S29i5[1];
			s29[mod*i+5+mod/2] <= _S29i5[0];
			s29[mod*i+6] <= _S29i6[1];
			s29[mod*i+6+mod/2] <= _S29i6[0];
			s29[mod*i+7] <= _S29i7[1];
			s29[mod*i+7+mod/2] <= _S29i7[0];
			s29[mod*i+8] <= _S29i8[1];
			s29[mod*i+8+mod/2] <= _S29i8[0];
			s29[mod*i+9] <= _S29i9[1];
			s29[mod*i+9+mod/2] <= _S29i9[0];
			s29[mod*i+10] <= _S29i10[1];
			s29[mod*i+10+mod/2] <= _S29i10[0];
			s29[mod*i+11] <= _S29i11[1];
			s29[mod*i+11+mod/2] <= _S29i11[0];
			s29[mod*i+12] <= _S29i12[1];
			s29[mod*i+12+mod/2] <= _S29i12[0];
			s29[mod*i+13] <= _S29i13[1];
			s29[mod*i+13+mod/2] <= _S29i13[0];
			s29[mod*i+14] <= _S29i14[1];
			s29[mod*i+14+mod/2] <= _S29i14[0];
			s29[mod*i+15] <= _S29i15[1];
			s29[mod*i+15+mod/2] <= _S29i15[0];
			s29[mod*i+16] <= _S29i16[1];
			s29[mod*i+16+mod/2] <= _S29i16[0];
			s29[mod*i+17] <= _S29i17[1];
			s29[mod*i+17+mod/2] <= _S29i17[0];
			s29[mod*i+18] <= _S29i18[1];
			s29[mod*i+18+mod/2] <= _S29i18[0];
			s29[mod*i+19] <= _S29i19[1];
			s29[mod*i+19+mod/2] <= _S29i19[0];
			s29[mod*i+20] <= _S29i20[1];
			s29[mod*i+20+mod/2] <= _S29i20[0];
			s29[mod*i+21] <= _S29i21[1];
			s29[mod*i+21+mod/2] <= _S29i21[0];
			s29[mod*i+22] <= _S29i22[1];
			s29[mod*i+22+mod/2] <= _S29i22[0];
			s29[mod*i+23] <= _S29i23[1];
			s29[mod*i+23+mod/2] <= _S29i23[0];
			s29[mod*i+24] <= _S29i24[1];
			s29[mod*i+24+mod/2] <= _S29i24[0];
			s29[mod*i+25] <= _S29i25[1];
			s29[mod*i+25+mod/2] <= _S29i25[0];
			s29[mod*i+26] <= _S29i26[1];
			s29[mod*i+26+mod/2] <= _S29i26[0];
			s29[mod*i+27] <= _S29i27[1];
			s29[mod*i+27+mod/2] <= _S29i27[0];
			s29[mod*i+28] <= _S29i28[1];
			s29[mod*i+28+mod/2] <= _S29i28[0];
			s29[mod*i+29] <= _S29i29[1];
			s29[mod*i+29+mod/2] <= _S29i29[0];
			s29[mod*i+30] <= _S29i30[1];
			s29[mod*i+30+mod/2] <= _S29i30[0];
			s29[mod*i+31] <= _S29i31[1];
			s29[mod*i+31+mod/2] <= _S29i31[0];
			s29[mod*i+32] <= _S29i32[1];
			s29[mod*i+32+mod/2] <= _S29i32[0];
			s29[mod*i+33] <= _S29i33[1];
			s29[mod*i+33+mod/2] <= _S29i33[0];
			s29[mod*i+34] <= _S29i34[1];
			s29[mod*i+34+mod/2] <= _S29i34[0];
			s29[mod*i+35] <= _S29i35[1];
			s29[mod*i+35+mod/2] <= _S29i35[0];
			s29[mod*i+36] <= _S29i36[1];
			s29[mod*i+36+mod/2] <= _S29i36[0];
			s29[mod*i+37] <= _S29i37[1];
			s29[mod*i+37+mod/2] <= _S29i37[0];
			s29[mod*i+38] <= _S29i38[1];
			s29[mod*i+38+mod/2] <= _S29i38[0];
			s29[mod*i+39] <= _S29i39[1];
			s29[mod*i+39+mod/2] <= _S29i39[0];
			s29[mod*i+40] <= _S29i40[1];
			s29[mod*i+40+mod/2] <= _S29i40[0];
			s29[mod*i+41] <= _S29i41[1];
			s29[mod*i+41+mod/2] <= _S29i41[0];
			s29[mod*i+42] <= _S29i42[1];
			s29[mod*i+42+mod/2] <= _S29i42[0];
			s29[mod*i+43] <= _S29i43[1];
			s29[mod*i+43+mod/2] <= _S29i43[0];
			s29[mod*i+44] <= _S29i44[1];
			s29[mod*i+44+mod/2] <= _S29i44[0];
			s29[mod*i+45] <= _S29i45[1];
			s29[mod*i+45+mod/2] <= _S29i45[0];
			s29[mod*i+46] <= _S29i46[1];
			s29[mod*i+46+mod/2] <= _S29i46[0];
			s29[mod*i+47] <= _S29i47[1];
			s29[mod*i+47+mod/2] <= _S29i47[0];
			s29[mod*i+48] <= _S29i48[1];
			s29[mod*i+48+mod/2] <= _S29i48[0];
			s29[mod*i+49] <= _S29i49[1];
			s29[mod*i+49+mod/2] <= _S29i49[0];
			s29[mod*i+50] <= _S29i50[1];
			s29[mod*i+50+mod/2] <= _S29i50[0];
			s29[mod*i+51] <= _S29i51[1];
			s29[mod*i+51+mod/2] <= _S29i51[0];
			s29[mod*i+52] <= _S29i52[1];
			s29[mod*i+52+mod/2] <= _S29i52[0];
			s29[mod*i+53] <= _S29i53[1];
			s29[mod*i+53+mod/2] <= _S29i53[0];
			s29[mod*i+54] <= _S29i54[1];
			s29[mod*i+54+mod/2] <= _S29i54[0];
			s29[mod*i+55] <= _S29i55[1];
			s29[mod*i+55+mod/2] <= _S29i55[0];
			s29[mod*i+56] <= _S29i56[1];
			s29[mod*i+56+mod/2] <= _S29i56[0];
			s29[mod*i+57] <= _S29i57[1];
			s29[mod*i+57+mod/2] <= _S29i57[0];
			s29[mod*i+58] <= _S29i58[1];
			s29[mod*i+58+mod/2] <= _S29i58[0];
			s29[mod*i+59] <= _S29i59[1];
			s29[mod*i+59+mod/2] <= _S29i59[0];
			s29[mod*i+60] <= _S29i60[1];
			s29[mod*i+60+mod/2] <= _S29i60[0];
			s29[mod*i+61] <= _S29i61[1];
			s29[mod*i+61+mod/2] <= _S29i61[0];
			s29[mod*i+62] <= _S29i62[1];
			s29[mod*i+62+mod/2] <= _S29i62[0];
			s29[mod*i+63] <= _S29i63[1];
			s29[mod*i+63+mod/2] <= _S29i63[0];
			s29[mod*i+64] <= _S29i64[1];
			s29[mod*i+64+mod/2] <= _S29i64[0];
			s29[mod*i+65] <= _S29i65[1];
			s29[mod*i+65+mod/2] <= _S29i65[0];
			s29[mod*i+66] <= _S29i66[1];
			s29[mod*i+66+mod/2] <= _S29i66[0];
			s29[mod*i+67] <= _S29i67[1];
			s29[mod*i+67+mod/2] <= _S29i67[0];
			s29[mod*i+68] <= _S29i68[1];
			s29[mod*i+68+mod/2] <= _S29i68[0];
			s29[mod*i+69] <= _S29i69[1];
			s29[mod*i+69+mod/2] <= _S29i69[0];
			s29[mod*i+70] <= _S29i70[1];
			s29[mod*i+70+mod/2] <= _S29i70[0];
			s29[mod*i+71] <= _S29i71[1];
			s29[mod*i+71+mod/2] <= _S29i71[0];
			s29[mod*i+72] <= _S29i72[1];
			s29[mod*i+72+mod/2] <= _S29i72[0];
			s29[mod*i+73] <= _S29i73[1];
			s29[mod*i+73+mod/2] <= _S29i73[0];
			s29[mod*i+74] <= _S29i74[1];
			s29[mod*i+74+mod/2] <= _S29i74[0];
			s29[mod*i+75] <= _S29i75[1];
			s29[mod*i+75+mod/2] <= _S29i75[0];
			s29[mod*i+76] <= _S29i76[1];
			s29[mod*i+76+mod/2] <= _S29i76[0];
			s29[mod*i+77] <= _S29i77[1];
			s29[mod*i+77+mod/2] <= _S29i77[0];
			s29[mod*i+78] <= _S29i78[1];
			s29[mod*i+78+mod/2] <= _S29i78[0];
			s29[mod*i+79] <= _S29i79[1];
			s29[mod*i+79+mod/2] <= _S29i79[0];
			s29[mod*i+80] <= _S29i80[1];
			s29[mod*i+80+mod/2] <= _S29i80[0];
			s29[mod*i+81] <= _S29i81[1];
			s29[mod*i+81+mod/2] <= _S29i81[0];
			s29[mod*i+82] <= _S29i82[1];
			s29[mod*i+82+mod/2] <= _S29i82[0];
			s29[mod*i+83] <= _S29i83[1];
			s29[mod*i+83+mod/2] <= _S29i83[0];
			s29[mod*i+84] <= _S29i84[1];
			s29[mod*i+84+mod/2] <= _S29i84[0];
			s29[mod*i+85] <= _S29i85[1];
			s29[mod*i+85+mod/2] <= _S29i85[0];
			s29[mod*i+86] <= _S29i86[1];
			s29[mod*i+86+mod/2] <= _S29i86[0];
			s29[mod*i+87] <= _S29i87[1];
			s29[mod*i+87+mod/2] <= _S29i87[0];
			s29[mod*i+88] <= _S29i88[1];
			s29[mod*i+88+mod/2] <= _S29i88[0];
			s29[mod*i+89] <= _S29i89[1];
			s29[mod*i+89+mod/2] <= _S29i89[0];
			s29[mod*i+90] <= _S29i90[1];
			s29[mod*i+90+mod/2] <= _S29i90[0];
			s29[mod*i+91] <= _S29i91[1];
			s29[mod*i+91+mod/2] <= _S29i91[0];
			s29[mod*i+92] <= _S29i92[1];
			s29[mod*i+92+mod/2] <= _S29i92[0];
			s29[mod*i+93] <= _S29i93[1];
			s29[mod*i+93+mod/2] <= _S29i93[0];
			s29[mod*i+94] <= _S29i94[1];
			s29[mod*i+94+mod/2] <= _S29i94[0];
			s29[mod*i+95] <= _S29i95[1];
			s29[mod*i+95+mod/2] <= _S29i95[0];
			s29[mod*i+96] <= _S29i96[1];
			s29[mod*i+96+mod/2] <= _S29i96[0];
			s29[mod*i+97] <= _S29i97[1];
			s29[mod*i+97+mod/2] <= _S29i97[0];
			s29[mod*i+98] <= _S29i98[1];
			s29[mod*i+98+mod/2] <= _S29i98[0];
			s29[mod*i+99] <= _S29i99[1];
			s29[mod*i+99+mod/2] <= _S29i99[0];
			s29[mod*i+100] <= _S29i100[1];
			s29[mod*i+100+mod/2] <= _S29i100[0];
			s29[mod*i+101] <= _S29i101[1];
			s29[mod*i+101+mod/2] <= _S29i101[0];
			s29[mod*i+102] <= _S29i102[1];
			s29[mod*i+102+mod/2] <= _S29i102[0];
			s29[mod*i+103] <= _S29i103[1];
			s29[mod*i+103+mod/2] <= _S29i103[0];
			s29[mod*i+104] <= _S29i104[1];
			s29[mod*i+104+mod/2] <= _S29i104[0];
			s29[mod*i+105] <= _S29i105[1];
			s29[mod*i+105+mod/2] <= _S29i105[0];
			s29[mod*i+106] <= _S29i106[1];
			s29[mod*i+106+mod/2] <= _S29i106[0];
			s29[mod*i+107] <= _S29i107[1];
			s29[mod*i+107+mod/2] <= _S29i107[0];
			s29[mod*i+108] <= _S29i108[1];
			s29[mod*i+108+mod/2] <= _S29i108[0];
			s29[mod*i+109] <= _S29i109[1];
			s29[mod*i+109+mod/2] <= _S29i109[0];
			s29[mod*i+110] <= _S29i110[1];
			s29[mod*i+110+mod/2] <= _S29i110[0];
			s29[mod*i+111] <= _S29i111[1];
			s29[mod*i+111+mod/2] <= _S29i111[0];
			s29[mod*i+112] <= _S29i112[1];
			s29[mod*i+112+mod/2] <= _S29i112[0];
			s29[mod*i+113] <= _S29i113[1];
			s29[mod*i+113+mod/2] <= _S29i113[0];
			s29[mod*i+114] <= _S29i114[1];
			s29[mod*i+114+mod/2] <= _S29i114[0];
			s29[mod*i+115] <= _S29i115[1];
			s29[mod*i+115+mod/2] <= _S29i115[0];
			s29[mod*i+116] <= _S29i116[1];
			s29[mod*i+116+mod/2] <= _S29i116[0];
			s29[mod*i+117] <= _S29i117[1];
			s29[mod*i+117+mod/2] <= _S29i117[0];
			s29[mod*i+118] <= _S29i118[1];
			s29[mod*i+118+mod/2] <= _S29i118[0];
			s29[mod*i+119] <= _S29i119[1];
			s29[mod*i+119+mod/2] <= _S29i119[0];
			s29[mod*i+120] <= _S29i120[1];
			s29[mod*i+120+mod/2] <= _S29i120[0];
			s29[mod*i+121] <= _S29i121[1];
			s29[mod*i+121+mod/2] <= _S29i121[0];
			s29[mod*i+122] <= _S29i122[1];
			s29[mod*i+122+mod/2] <= _S29i122[0];
			s29[mod*i+123] <= _S29i123[1];
			s29[mod*i+123+mod/2] <= _S29i123[0];
			s29[mod*i+124] <= _S29i124[1];
			s29[mod*i+124+mod/2] <= _S29i124[0];
			s29[mod*i+125] <= _S29i125[1];
			s29[mod*i+125+mod/2] <= _S29i125[0];
			s29[mod*i+126] <= _S29i126[1];
			s29[mod*i+126+mod/2] <= _S29i126[0];
			s29[mod*i+127] <= _S29i127[1];
			s29[mod*i+127+mod/2] <= _S29i127[0];
		end
	end
	p29.enq(1);
endrule
rule _Q77;
	p29.deq;
	let mod = 128;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S30i0 = min_max(pack(s29[mod*i+0]) , pack(s29[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S30i1 = min_max(pack(s29[mod*i+1]) , pack(s29[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S30i2 = min_max(pack(s29[mod*i+2]) , pack(s29[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S30i3 = min_max(pack(s29[mod*i+3]) , pack(s29[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S30i4 = min_max(pack(s29[mod*i+4]) , pack(s29[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S30i5 = min_max(pack(s29[mod*i+5]) , pack(s29[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S30i6 = min_max(pack(s29[mod*i+6]) , pack(s29[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S30i7 = min_max(pack(s29[mod*i+7]) , pack(s29[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S30i8 = min_max(pack(s29[mod*i+8]) , pack(s29[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S30i9 = min_max(pack(s29[mod*i+9]) , pack(s29[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S30i10 = min_max(pack(s29[mod*i+10]) , pack(s29[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S30i11 = min_max(pack(s29[mod*i+11]) , pack(s29[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S30i12 = min_max(pack(s29[mod*i+12]) , pack(s29[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S30i13 = min_max(pack(s29[mod*i+13]) , pack(s29[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S30i14 = min_max(pack(s29[mod*i+14]) , pack(s29[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S30i15 = min_max(pack(s29[mod*i+15]) , pack(s29[mod*i+15+mod/2]));
			 Vector#(2, Int#(32)) _S30i16 = min_max(pack(s29[mod*i+16]) , pack(s29[mod*i+16+mod/2]));
			 Vector#(2, Int#(32)) _S30i17 = min_max(pack(s29[mod*i+17]) , pack(s29[mod*i+17+mod/2]));
			 Vector#(2, Int#(32)) _S30i18 = min_max(pack(s29[mod*i+18]) , pack(s29[mod*i+18+mod/2]));
			 Vector#(2, Int#(32)) _S30i19 = min_max(pack(s29[mod*i+19]) , pack(s29[mod*i+19+mod/2]));
			 Vector#(2, Int#(32)) _S30i20 = min_max(pack(s29[mod*i+20]) , pack(s29[mod*i+20+mod/2]));
			 Vector#(2, Int#(32)) _S30i21 = min_max(pack(s29[mod*i+21]) , pack(s29[mod*i+21+mod/2]));
			 Vector#(2, Int#(32)) _S30i22 = min_max(pack(s29[mod*i+22]) , pack(s29[mod*i+22+mod/2]));
			 Vector#(2, Int#(32)) _S30i23 = min_max(pack(s29[mod*i+23]) , pack(s29[mod*i+23+mod/2]));
			 Vector#(2, Int#(32)) _S30i24 = min_max(pack(s29[mod*i+24]) , pack(s29[mod*i+24+mod/2]));
			 Vector#(2, Int#(32)) _S30i25 = min_max(pack(s29[mod*i+25]) , pack(s29[mod*i+25+mod/2]));
			 Vector#(2, Int#(32)) _S30i26 = min_max(pack(s29[mod*i+26]) , pack(s29[mod*i+26+mod/2]));
			 Vector#(2, Int#(32)) _S30i27 = min_max(pack(s29[mod*i+27]) , pack(s29[mod*i+27+mod/2]));
			 Vector#(2, Int#(32)) _S30i28 = min_max(pack(s29[mod*i+28]) , pack(s29[mod*i+28+mod/2]));
			 Vector#(2, Int#(32)) _S30i29 = min_max(pack(s29[mod*i+29]) , pack(s29[mod*i+29+mod/2]));
			 Vector#(2, Int#(32)) _S30i30 = min_max(pack(s29[mod*i+30]) , pack(s29[mod*i+30+mod/2]));
			 Vector#(2, Int#(32)) _S30i31 = min_max(pack(s29[mod*i+31]) , pack(s29[mod*i+31+mod/2]));
			 Vector#(2, Int#(32)) _S30i32 = min_max(pack(s29[mod*i+32]) , pack(s29[mod*i+32+mod/2]));
			 Vector#(2, Int#(32)) _S30i33 = min_max(pack(s29[mod*i+33]) , pack(s29[mod*i+33+mod/2]));
			 Vector#(2, Int#(32)) _S30i34 = min_max(pack(s29[mod*i+34]) , pack(s29[mod*i+34+mod/2]));
			 Vector#(2, Int#(32)) _S30i35 = min_max(pack(s29[mod*i+35]) , pack(s29[mod*i+35+mod/2]));
			 Vector#(2, Int#(32)) _S30i36 = min_max(pack(s29[mod*i+36]) , pack(s29[mod*i+36+mod/2]));
			 Vector#(2, Int#(32)) _S30i37 = min_max(pack(s29[mod*i+37]) , pack(s29[mod*i+37+mod/2]));
			 Vector#(2, Int#(32)) _S30i38 = min_max(pack(s29[mod*i+38]) , pack(s29[mod*i+38+mod/2]));
			 Vector#(2, Int#(32)) _S30i39 = min_max(pack(s29[mod*i+39]) , pack(s29[mod*i+39+mod/2]));
			 Vector#(2, Int#(32)) _S30i40 = min_max(pack(s29[mod*i+40]) , pack(s29[mod*i+40+mod/2]));
			 Vector#(2, Int#(32)) _S30i41 = min_max(pack(s29[mod*i+41]) , pack(s29[mod*i+41+mod/2]));
			 Vector#(2, Int#(32)) _S30i42 = min_max(pack(s29[mod*i+42]) , pack(s29[mod*i+42+mod/2]));
			 Vector#(2, Int#(32)) _S30i43 = min_max(pack(s29[mod*i+43]) , pack(s29[mod*i+43+mod/2]));
			 Vector#(2, Int#(32)) _S30i44 = min_max(pack(s29[mod*i+44]) , pack(s29[mod*i+44+mod/2]));
			 Vector#(2, Int#(32)) _S30i45 = min_max(pack(s29[mod*i+45]) , pack(s29[mod*i+45+mod/2]));
			 Vector#(2, Int#(32)) _S30i46 = min_max(pack(s29[mod*i+46]) , pack(s29[mod*i+46+mod/2]));
			 Vector#(2, Int#(32)) _S30i47 = min_max(pack(s29[mod*i+47]) , pack(s29[mod*i+47+mod/2]));
			 Vector#(2, Int#(32)) _S30i48 = min_max(pack(s29[mod*i+48]) , pack(s29[mod*i+48+mod/2]));
			 Vector#(2, Int#(32)) _S30i49 = min_max(pack(s29[mod*i+49]) , pack(s29[mod*i+49+mod/2]));
			 Vector#(2, Int#(32)) _S30i50 = min_max(pack(s29[mod*i+50]) , pack(s29[mod*i+50+mod/2]));
			 Vector#(2, Int#(32)) _S30i51 = min_max(pack(s29[mod*i+51]) , pack(s29[mod*i+51+mod/2]));
			 Vector#(2, Int#(32)) _S30i52 = min_max(pack(s29[mod*i+52]) , pack(s29[mod*i+52+mod/2]));
			 Vector#(2, Int#(32)) _S30i53 = min_max(pack(s29[mod*i+53]) , pack(s29[mod*i+53+mod/2]));
			 Vector#(2, Int#(32)) _S30i54 = min_max(pack(s29[mod*i+54]) , pack(s29[mod*i+54+mod/2]));
			 Vector#(2, Int#(32)) _S30i55 = min_max(pack(s29[mod*i+55]) , pack(s29[mod*i+55+mod/2]));
			 Vector#(2, Int#(32)) _S30i56 = min_max(pack(s29[mod*i+56]) , pack(s29[mod*i+56+mod/2]));
			 Vector#(2, Int#(32)) _S30i57 = min_max(pack(s29[mod*i+57]) , pack(s29[mod*i+57+mod/2]));
			 Vector#(2, Int#(32)) _S30i58 = min_max(pack(s29[mod*i+58]) , pack(s29[mod*i+58+mod/2]));
			 Vector#(2, Int#(32)) _S30i59 = min_max(pack(s29[mod*i+59]) , pack(s29[mod*i+59+mod/2]));
			 Vector#(2, Int#(32)) _S30i60 = min_max(pack(s29[mod*i+60]) , pack(s29[mod*i+60+mod/2]));
			 Vector#(2, Int#(32)) _S30i61 = min_max(pack(s29[mod*i+61]) , pack(s29[mod*i+61+mod/2]));
			 Vector#(2, Int#(32)) _S30i62 = min_max(pack(s29[mod*i+62]) , pack(s29[mod*i+62+mod/2]));
			 Vector#(2, Int#(32)) _S30i63 = min_max(pack(s29[mod*i+63]) , pack(s29[mod*i+63+mod/2]));
		if ((i/2)%2 == 0) begin
			s30[mod*i+0] <= _S30i0[0];
			s30[mod*i+0+mod/2] <= _S30i0[1];
			s30[mod*i+1] <= _S30i1[0];
			s30[mod*i+1+mod/2] <= _S30i1[1];
			s30[mod*i+2] <= _S30i2[0];
			s30[mod*i+2+mod/2] <= _S30i2[1];
			s30[mod*i+3] <= _S30i3[0];
			s30[mod*i+3+mod/2] <= _S30i3[1];
			s30[mod*i+4] <= _S30i4[0];
			s30[mod*i+4+mod/2] <= _S30i4[1];
			s30[mod*i+5] <= _S30i5[0];
			s30[mod*i+5+mod/2] <= _S30i5[1];
			s30[mod*i+6] <= _S30i6[0];
			s30[mod*i+6+mod/2] <= _S30i6[1];
			s30[mod*i+7] <= _S30i7[0];
			s30[mod*i+7+mod/2] <= _S30i7[1];
			s30[mod*i+8] <= _S30i8[0];
			s30[mod*i+8+mod/2] <= _S30i8[1];
			s30[mod*i+9] <= _S30i9[0];
			s30[mod*i+9+mod/2] <= _S30i9[1];
			s30[mod*i+10] <= _S30i10[0];
			s30[mod*i+10+mod/2] <= _S30i10[1];
			s30[mod*i+11] <= _S30i11[0];
			s30[mod*i+11+mod/2] <= _S30i11[1];
			s30[mod*i+12] <= _S30i12[0];
			s30[mod*i+12+mod/2] <= _S30i12[1];
			s30[mod*i+13] <= _S30i13[0];
			s30[mod*i+13+mod/2] <= _S30i13[1];
			s30[mod*i+14] <= _S30i14[0];
			s30[mod*i+14+mod/2] <= _S30i14[1];
			s30[mod*i+15] <= _S30i15[0];
			s30[mod*i+15+mod/2] <= _S30i15[1];
			s30[mod*i+16] <= _S30i16[0];
			s30[mod*i+16+mod/2] <= _S30i16[1];
			s30[mod*i+17] <= _S30i17[0];
			s30[mod*i+17+mod/2] <= _S30i17[1];
			s30[mod*i+18] <= _S30i18[0];
			s30[mod*i+18+mod/2] <= _S30i18[1];
			s30[mod*i+19] <= _S30i19[0];
			s30[mod*i+19+mod/2] <= _S30i19[1];
			s30[mod*i+20] <= _S30i20[0];
			s30[mod*i+20+mod/2] <= _S30i20[1];
			s30[mod*i+21] <= _S30i21[0];
			s30[mod*i+21+mod/2] <= _S30i21[1];
			s30[mod*i+22] <= _S30i22[0];
			s30[mod*i+22+mod/2] <= _S30i22[1];
			s30[mod*i+23] <= _S30i23[0];
			s30[mod*i+23+mod/2] <= _S30i23[1];
			s30[mod*i+24] <= _S30i24[0];
			s30[mod*i+24+mod/2] <= _S30i24[1];
			s30[mod*i+25] <= _S30i25[0];
			s30[mod*i+25+mod/2] <= _S30i25[1];
			s30[mod*i+26] <= _S30i26[0];
			s30[mod*i+26+mod/2] <= _S30i26[1];
			s30[mod*i+27] <= _S30i27[0];
			s30[mod*i+27+mod/2] <= _S30i27[1];
			s30[mod*i+28] <= _S30i28[0];
			s30[mod*i+28+mod/2] <= _S30i28[1];
			s30[mod*i+29] <= _S30i29[0];
			s30[mod*i+29+mod/2] <= _S30i29[1];
			s30[mod*i+30] <= _S30i30[0];
			s30[mod*i+30+mod/2] <= _S30i30[1];
			s30[mod*i+31] <= _S30i31[0];
			s30[mod*i+31+mod/2] <= _S30i31[1];
			s30[mod*i+32] <= _S30i32[0];
			s30[mod*i+32+mod/2] <= _S30i32[1];
			s30[mod*i+33] <= _S30i33[0];
			s30[mod*i+33+mod/2] <= _S30i33[1];
			s30[mod*i+34] <= _S30i34[0];
			s30[mod*i+34+mod/2] <= _S30i34[1];
			s30[mod*i+35] <= _S30i35[0];
			s30[mod*i+35+mod/2] <= _S30i35[1];
			s30[mod*i+36] <= _S30i36[0];
			s30[mod*i+36+mod/2] <= _S30i36[1];
			s30[mod*i+37] <= _S30i37[0];
			s30[mod*i+37+mod/2] <= _S30i37[1];
			s30[mod*i+38] <= _S30i38[0];
			s30[mod*i+38+mod/2] <= _S30i38[1];
			s30[mod*i+39] <= _S30i39[0];
			s30[mod*i+39+mod/2] <= _S30i39[1];
			s30[mod*i+40] <= _S30i40[0];
			s30[mod*i+40+mod/2] <= _S30i40[1];
			s30[mod*i+41] <= _S30i41[0];
			s30[mod*i+41+mod/2] <= _S30i41[1];
			s30[mod*i+42] <= _S30i42[0];
			s30[mod*i+42+mod/2] <= _S30i42[1];
			s30[mod*i+43] <= _S30i43[0];
			s30[mod*i+43+mod/2] <= _S30i43[1];
			s30[mod*i+44] <= _S30i44[0];
			s30[mod*i+44+mod/2] <= _S30i44[1];
			s30[mod*i+45] <= _S30i45[0];
			s30[mod*i+45+mod/2] <= _S30i45[1];
			s30[mod*i+46] <= _S30i46[0];
			s30[mod*i+46+mod/2] <= _S30i46[1];
			s30[mod*i+47] <= _S30i47[0];
			s30[mod*i+47+mod/2] <= _S30i47[1];
			s30[mod*i+48] <= _S30i48[0];
			s30[mod*i+48+mod/2] <= _S30i48[1];
			s30[mod*i+49] <= _S30i49[0];
			s30[mod*i+49+mod/2] <= _S30i49[1];
			s30[mod*i+50] <= _S30i50[0];
			s30[mod*i+50+mod/2] <= _S30i50[1];
			s30[mod*i+51] <= _S30i51[0];
			s30[mod*i+51+mod/2] <= _S30i51[1];
			s30[mod*i+52] <= _S30i52[0];
			s30[mod*i+52+mod/2] <= _S30i52[1];
			s30[mod*i+53] <= _S30i53[0];
			s30[mod*i+53+mod/2] <= _S30i53[1];
			s30[mod*i+54] <= _S30i54[0];
			s30[mod*i+54+mod/2] <= _S30i54[1];
			s30[mod*i+55] <= _S30i55[0];
			s30[mod*i+55+mod/2] <= _S30i55[1];
			s30[mod*i+56] <= _S30i56[0];
			s30[mod*i+56+mod/2] <= _S30i56[1];
			s30[mod*i+57] <= _S30i57[0];
			s30[mod*i+57+mod/2] <= _S30i57[1];
			s30[mod*i+58] <= _S30i58[0];
			s30[mod*i+58+mod/2] <= _S30i58[1];
			s30[mod*i+59] <= _S30i59[0];
			s30[mod*i+59+mod/2] <= _S30i59[1];
			s30[mod*i+60] <= _S30i60[0];
			s30[mod*i+60+mod/2] <= _S30i60[1];
			s30[mod*i+61] <= _S30i61[0];
			s30[mod*i+61+mod/2] <= _S30i61[1];
			s30[mod*i+62] <= _S30i62[0];
			s30[mod*i+62+mod/2] <= _S30i62[1];
			s30[mod*i+63] <= _S30i63[0];
			s30[mod*i+63+mod/2] <= _S30i63[1];
		end
		else begin
			s30[mod*i+0] <= _S30i0[1];
			s30[mod*i+0+mod/2] <= _S30i0[0];
			s30[mod*i+1] <= _S30i1[1];
			s30[mod*i+1+mod/2] <= _S30i1[0];
			s30[mod*i+2] <= _S30i2[1];
			s30[mod*i+2+mod/2] <= _S30i2[0];
			s30[mod*i+3] <= _S30i3[1];
			s30[mod*i+3+mod/2] <= _S30i3[0];
			s30[mod*i+4] <= _S30i4[1];
			s30[mod*i+4+mod/2] <= _S30i4[0];
			s30[mod*i+5] <= _S30i5[1];
			s30[mod*i+5+mod/2] <= _S30i5[0];
			s30[mod*i+6] <= _S30i6[1];
			s30[mod*i+6+mod/2] <= _S30i6[0];
			s30[mod*i+7] <= _S30i7[1];
			s30[mod*i+7+mod/2] <= _S30i7[0];
			s30[mod*i+8] <= _S30i8[1];
			s30[mod*i+8+mod/2] <= _S30i8[0];
			s30[mod*i+9] <= _S30i9[1];
			s30[mod*i+9+mod/2] <= _S30i9[0];
			s30[mod*i+10] <= _S30i10[1];
			s30[mod*i+10+mod/2] <= _S30i10[0];
			s30[mod*i+11] <= _S30i11[1];
			s30[mod*i+11+mod/2] <= _S30i11[0];
			s30[mod*i+12] <= _S30i12[1];
			s30[mod*i+12+mod/2] <= _S30i12[0];
			s30[mod*i+13] <= _S30i13[1];
			s30[mod*i+13+mod/2] <= _S30i13[0];
			s30[mod*i+14] <= _S30i14[1];
			s30[mod*i+14+mod/2] <= _S30i14[0];
			s30[mod*i+15] <= _S30i15[1];
			s30[mod*i+15+mod/2] <= _S30i15[0];
			s30[mod*i+16] <= _S30i16[1];
			s30[mod*i+16+mod/2] <= _S30i16[0];
			s30[mod*i+17] <= _S30i17[1];
			s30[mod*i+17+mod/2] <= _S30i17[0];
			s30[mod*i+18] <= _S30i18[1];
			s30[mod*i+18+mod/2] <= _S30i18[0];
			s30[mod*i+19] <= _S30i19[1];
			s30[mod*i+19+mod/2] <= _S30i19[0];
			s30[mod*i+20] <= _S30i20[1];
			s30[mod*i+20+mod/2] <= _S30i20[0];
			s30[mod*i+21] <= _S30i21[1];
			s30[mod*i+21+mod/2] <= _S30i21[0];
			s30[mod*i+22] <= _S30i22[1];
			s30[mod*i+22+mod/2] <= _S30i22[0];
			s30[mod*i+23] <= _S30i23[1];
			s30[mod*i+23+mod/2] <= _S30i23[0];
			s30[mod*i+24] <= _S30i24[1];
			s30[mod*i+24+mod/2] <= _S30i24[0];
			s30[mod*i+25] <= _S30i25[1];
			s30[mod*i+25+mod/2] <= _S30i25[0];
			s30[mod*i+26] <= _S30i26[1];
			s30[mod*i+26+mod/2] <= _S30i26[0];
			s30[mod*i+27] <= _S30i27[1];
			s30[mod*i+27+mod/2] <= _S30i27[0];
			s30[mod*i+28] <= _S30i28[1];
			s30[mod*i+28+mod/2] <= _S30i28[0];
			s30[mod*i+29] <= _S30i29[1];
			s30[mod*i+29+mod/2] <= _S30i29[0];
			s30[mod*i+30] <= _S30i30[1];
			s30[mod*i+30+mod/2] <= _S30i30[0];
			s30[mod*i+31] <= _S30i31[1];
			s30[mod*i+31+mod/2] <= _S30i31[0];
			s30[mod*i+32] <= _S30i32[1];
			s30[mod*i+32+mod/2] <= _S30i32[0];
			s30[mod*i+33] <= _S30i33[1];
			s30[mod*i+33+mod/2] <= _S30i33[0];
			s30[mod*i+34] <= _S30i34[1];
			s30[mod*i+34+mod/2] <= _S30i34[0];
			s30[mod*i+35] <= _S30i35[1];
			s30[mod*i+35+mod/2] <= _S30i35[0];
			s30[mod*i+36] <= _S30i36[1];
			s30[mod*i+36+mod/2] <= _S30i36[0];
			s30[mod*i+37] <= _S30i37[1];
			s30[mod*i+37+mod/2] <= _S30i37[0];
			s30[mod*i+38] <= _S30i38[1];
			s30[mod*i+38+mod/2] <= _S30i38[0];
			s30[mod*i+39] <= _S30i39[1];
			s30[mod*i+39+mod/2] <= _S30i39[0];
			s30[mod*i+40] <= _S30i40[1];
			s30[mod*i+40+mod/2] <= _S30i40[0];
			s30[mod*i+41] <= _S30i41[1];
			s30[mod*i+41+mod/2] <= _S30i41[0];
			s30[mod*i+42] <= _S30i42[1];
			s30[mod*i+42+mod/2] <= _S30i42[0];
			s30[mod*i+43] <= _S30i43[1];
			s30[mod*i+43+mod/2] <= _S30i43[0];
			s30[mod*i+44] <= _S30i44[1];
			s30[mod*i+44+mod/2] <= _S30i44[0];
			s30[mod*i+45] <= _S30i45[1];
			s30[mod*i+45+mod/2] <= _S30i45[0];
			s30[mod*i+46] <= _S30i46[1];
			s30[mod*i+46+mod/2] <= _S30i46[0];
			s30[mod*i+47] <= _S30i47[1];
			s30[mod*i+47+mod/2] <= _S30i47[0];
			s30[mod*i+48] <= _S30i48[1];
			s30[mod*i+48+mod/2] <= _S30i48[0];
			s30[mod*i+49] <= _S30i49[1];
			s30[mod*i+49+mod/2] <= _S30i49[0];
			s30[mod*i+50] <= _S30i50[1];
			s30[mod*i+50+mod/2] <= _S30i50[0];
			s30[mod*i+51] <= _S30i51[1];
			s30[mod*i+51+mod/2] <= _S30i51[0];
			s30[mod*i+52] <= _S30i52[1];
			s30[mod*i+52+mod/2] <= _S30i52[0];
			s30[mod*i+53] <= _S30i53[1];
			s30[mod*i+53+mod/2] <= _S30i53[0];
			s30[mod*i+54] <= _S30i54[1];
			s30[mod*i+54+mod/2] <= _S30i54[0];
			s30[mod*i+55] <= _S30i55[1];
			s30[mod*i+55+mod/2] <= _S30i55[0];
			s30[mod*i+56] <= _S30i56[1];
			s30[mod*i+56+mod/2] <= _S30i56[0];
			s30[mod*i+57] <= _S30i57[1];
			s30[mod*i+57+mod/2] <= _S30i57[0];
			s30[mod*i+58] <= _S30i58[1];
			s30[mod*i+58+mod/2] <= _S30i58[0];
			s30[mod*i+59] <= _S30i59[1];
			s30[mod*i+59+mod/2] <= _S30i59[0];
			s30[mod*i+60] <= _S30i60[1];
			s30[mod*i+60+mod/2] <= _S30i60[0];
			s30[mod*i+61] <= _S30i61[1];
			s30[mod*i+61+mod/2] <= _S30i61[0];
			s30[mod*i+62] <= _S30i62[1];
			s30[mod*i+62+mod/2] <= _S30i62[0];
			s30[mod*i+63] <= _S30i63[1];
			s30[mod*i+63+mod/2] <= _S30i63[0];
		end
	end
	p30.enq(1);
endrule
rule _Q76;
	p30.deq;
	let mod = 64;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S31i0 = min_max(pack(s30[mod*i+0]) , pack(s30[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S31i1 = min_max(pack(s30[mod*i+1]) , pack(s30[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S31i2 = min_max(pack(s30[mod*i+2]) , pack(s30[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S31i3 = min_max(pack(s30[mod*i+3]) , pack(s30[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S31i4 = min_max(pack(s30[mod*i+4]) , pack(s30[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S31i5 = min_max(pack(s30[mod*i+5]) , pack(s30[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S31i6 = min_max(pack(s30[mod*i+6]) , pack(s30[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S31i7 = min_max(pack(s30[mod*i+7]) , pack(s30[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S31i8 = min_max(pack(s30[mod*i+8]) , pack(s30[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S31i9 = min_max(pack(s30[mod*i+9]) , pack(s30[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S31i10 = min_max(pack(s30[mod*i+10]) , pack(s30[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S31i11 = min_max(pack(s30[mod*i+11]) , pack(s30[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S31i12 = min_max(pack(s30[mod*i+12]) , pack(s30[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S31i13 = min_max(pack(s30[mod*i+13]) , pack(s30[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S31i14 = min_max(pack(s30[mod*i+14]) , pack(s30[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S31i15 = min_max(pack(s30[mod*i+15]) , pack(s30[mod*i+15+mod/2]));
			 Vector#(2, Int#(32)) _S31i16 = min_max(pack(s30[mod*i+16]) , pack(s30[mod*i+16+mod/2]));
			 Vector#(2, Int#(32)) _S31i17 = min_max(pack(s30[mod*i+17]) , pack(s30[mod*i+17+mod/2]));
			 Vector#(2, Int#(32)) _S31i18 = min_max(pack(s30[mod*i+18]) , pack(s30[mod*i+18+mod/2]));
			 Vector#(2, Int#(32)) _S31i19 = min_max(pack(s30[mod*i+19]) , pack(s30[mod*i+19+mod/2]));
			 Vector#(2, Int#(32)) _S31i20 = min_max(pack(s30[mod*i+20]) , pack(s30[mod*i+20+mod/2]));
			 Vector#(2, Int#(32)) _S31i21 = min_max(pack(s30[mod*i+21]) , pack(s30[mod*i+21+mod/2]));
			 Vector#(2, Int#(32)) _S31i22 = min_max(pack(s30[mod*i+22]) , pack(s30[mod*i+22+mod/2]));
			 Vector#(2, Int#(32)) _S31i23 = min_max(pack(s30[mod*i+23]) , pack(s30[mod*i+23+mod/2]));
			 Vector#(2, Int#(32)) _S31i24 = min_max(pack(s30[mod*i+24]) , pack(s30[mod*i+24+mod/2]));
			 Vector#(2, Int#(32)) _S31i25 = min_max(pack(s30[mod*i+25]) , pack(s30[mod*i+25+mod/2]));
			 Vector#(2, Int#(32)) _S31i26 = min_max(pack(s30[mod*i+26]) , pack(s30[mod*i+26+mod/2]));
			 Vector#(2, Int#(32)) _S31i27 = min_max(pack(s30[mod*i+27]) , pack(s30[mod*i+27+mod/2]));
			 Vector#(2, Int#(32)) _S31i28 = min_max(pack(s30[mod*i+28]) , pack(s30[mod*i+28+mod/2]));
			 Vector#(2, Int#(32)) _S31i29 = min_max(pack(s30[mod*i+29]) , pack(s30[mod*i+29+mod/2]));
			 Vector#(2, Int#(32)) _S31i30 = min_max(pack(s30[mod*i+30]) , pack(s30[mod*i+30+mod/2]));
			 Vector#(2, Int#(32)) _S31i31 = min_max(pack(s30[mod*i+31]) , pack(s30[mod*i+31+mod/2]));
		if ((i/4)%2 == 0) begin
			s31[mod*i+0] <= _S31i0[0];
			s31[mod*i+0+mod/2] <= _S31i0[1];
			s31[mod*i+1] <= _S31i1[0];
			s31[mod*i+1+mod/2] <= _S31i1[1];
			s31[mod*i+2] <= _S31i2[0];
			s31[mod*i+2+mod/2] <= _S31i2[1];
			s31[mod*i+3] <= _S31i3[0];
			s31[mod*i+3+mod/2] <= _S31i3[1];
			s31[mod*i+4] <= _S31i4[0];
			s31[mod*i+4+mod/2] <= _S31i4[1];
			s31[mod*i+5] <= _S31i5[0];
			s31[mod*i+5+mod/2] <= _S31i5[1];
			s31[mod*i+6] <= _S31i6[0];
			s31[mod*i+6+mod/2] <= _S31i6[1];
			s31[mod*i+7] <= _S31i7[0];
			s31[mod*i+7+mod/2] <= _S31i7[1];
			s31[mod*i+8] <= _S31i8[0];
			s31[mod*i+8+mod/2] <= _S31i8[1];
			s31[mod*i+9] <= _S31i9[0];
			s31[mod*i+9+mod/2] <= _S31i9[1];
			s31[mod*i+10] <= _S31i10[0];
			s31[mod*i+10+mod/2] <= _S31i10[1];
			s31[mod*i+11] <= _S31i11[0];
			s31[mod*i+11+mod/2] <= _S31i11[1];
			s31[mod*i+12] <= _S31i12[0];
			s31[mod*i+12+mod/2] <= _S31i12[1];
			s31[mod*i+13] <= _S31i13[0];
			s31[mod*i+13+mod/2] <= _S31i13[1];
			s31[mod*i+14] <= _S31i14[0];
			s31[mod*i+14+mod/2] <= _S31i14[1];
			s31[mod*i+15] <= _S31i15[0];
			s31[mod*i+15+mod/2] <= _S31i15[1];
			s31[mod*i+16] <= _S31i16[0];
			s31[mod*i+16+mod/2] <= _S31i16[1];
			s31[mod*i+17] <= _S31i17[0];
			s31[mod*i+17+mod/2] <= _S31i17[1];
			s31[mod*i+18] <= _S31i18[0];
			s31[mod*i+18+mod/2] <= _S31i18[1];
			s31[mod*i+19] <= _S31i19[0];
			s31[mod*i+19+mod/2] <= _S31i19[1];
			s31[mod*i+20] <= _S31i20[0];
			s31[mod*i+20+mod/2] <= _S31i20[1];
			s31[mod*i+21] <= _S31i21[0];
			s31[mod*i+21+mod/2] <= _S31i21[1];
			s31[mod*i+22] <= _S31i22[0];
			s31[mod*i+22+mod/2] <= _S31i22[1];
			s31[mod*i+23] <= _S31i23[0];
			s31[mod*i+23+mod/2] <= _S31i23[1];
			s31[mod*i+24] <= _S31i24[0];
			s31[mod*i+24+mod/2] <= _S31i24[1];
			s31[mod*i+25] <= _S31i25[0];
			s31[mod*i+25+mod/2] <= _S31i25[1];
			s31[mod*i+26] <= _S31i26[0];
			s31[mod*i+26+mod/2] <= _S31i26[1];
			s31[mod*i+27] <= _S31i27[0];
			s31[mod*i+27+mod/2] <= _S31i27[1];
			s31[mod*i+28] <= _S31i28[0];
			s31[mod*i+28+mod/2] <= _S31i28[1];
			s31[mod*i+29] <= _S31i29[0];
			s31[mod*i+29+mod/2] <= _S31i29[1];
			s31[mod*i+30] <= _S31i30[0];
			s31[mod*i+30+mod/2] <= _S31i30[1];
			s31[mod*i+31] <= _S31i31[0];
			s31[mod*i+31+mod/2] <= _S31i31[1];
		end
		else begin
			s31[mod*i+0] <= _S31i0[1];
			s31[mod*i+0+mod/2] <= _S31i0[0];
			s31[mod*i+1] <= _S31i1[1];
			s31[mod*i+1+mod/2] <= _S31i1[0];
			s31[mod*i+2] <= _S31i2[1];
			s31[mod*i+2+mod/2] <= _S31i2[0];
			s31[mod*i+3] <= _S31i3[1];
			s31[mod*i+3+mod/2] <= _S31i3[0];
			s31[mod*i+4] <= _S31i4[1];
			s31[mod*i+4+mod/2] <= _S31i4[0];
			s31[mod*i+5] <= _S31i5[1];
			s31[mod*i+5+mod/2] <= _S31i5[0];
			s31[mod*i+6] <= _S31i6[1];
			s31[mod*i+6+mod/2] <= _S31i6[0];
			s31[mod*i+7] <= _S31i7[1];
			s31[mod*i+7+mod/2] <= _S31i7[0];
			s31[mod*i+8] <= _S31i8[1];
			s31[mod*i+8+mod/2] <= _S31i8[0];
			s31[mod*i+9] <= _S31i9[1];
			s31[mod*i+9+mod/2] <= _S31i9[0];
			s31[mod*i+10] <= _S31i10[1];
			s31[mod*i+10+mod/2] <= _S31i10[0];
			s31[mod*i+11] <= _S31i11[1];
			s31[mod*i+11+mod/2] <= _S31i11[0];
			s31[mod*i+12] <= _S31i12[1];
			s31[mod*i+12+mod/2] <= _S31i12[0];
			s31[mod*i+13] <= _S31i13[1];
			s31[mod*i+13+mod/2] <= _S31i13[0];
			s31[mod*i+14] <= _S31i14[1];
			s31[mod*i+14+mod/2] <= _S31i14[0];
			s31[mod*i+15] <= _S31i15[1];
			s31[mod*i+15+mod/2] <= _S31i15[0];
			s31[mod*i+16] <= _S31i16[1];
			s31[mod*i+16+mod/2] <= _S31i16[0];
			s31[mod*i+17] <= _S31i17[1];
			s31[mod*i+17+mod/2] <= _S31i17[0];
			s31[mod*i+18] <= _S31i18[1];
			s31[mod*i+18+mod/2] <= _S31i18[0];
			s31[mod*i+19] <= _S31i19[1];
			s31[mod*i+19+mod/2] <= _S31i19[0];
			s31[mod*i+20] <= _S31i20[1];
			s31[mod*i+20+mod/2] <= _S31i20[0];
			s31[mod*i+21] <= _S31i21[1];
			s31[mod*i+21+mod/2] <= _S31i21[0];
			s31[mod*i+22] <= _S31i22[1];
			s31[mod*i+22+mod/2] <= _S31i22[0];
			s31[mod*i+23] <= _S31i23[1];
			s31[mod*i+23+mod/2] <= _S31i23[0];
			s31[mod*i+24] <= _S31i24[1];
			s31[mod*i+24+mod/2] <= _S31i24[0];
			s31[mod*i+25] <= _S31i25[1];
			s31[mod*i+25+mod/2] <= _S31i25[0];
			s31[mod*i+26] <= _S31i26[1];
			s31[mod*i+26+mod/2] <= _S31i26[0];
			s31[mod*i+27] <= _S31i27[1];
			s31[mod*i+27+mod/2] <= _S31i27[0];
			s31[mod*i+28] <= _S31i28[1];
			s31[mod*i+28+mod/2] <= _S31i28[0];
			s31[mod*i+29] <= _S31i29[1];
			s31[mod*i+29+mod/2] <= _S31i29[0];
			s31[mod*i+30] <= _S31i30[1];
			s31[mod*i+30+mod/2] <= _S31i30[0];
			s31[mod*i+31] <= _S31i31[1];
			s31[mod*i+31+mod/2] <= _S31i31[0];
		end
	end
	p31.enq(1);
endrule
rule _Q75;
	p31.deq;
	let mod = 32;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S32i0 = min_max(pack(s31[mod*i+0]) , pack(s31[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S32i1 = min_max(pack(s31[mod*i+1]) , pack(s31[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S32i2 = min_max(pack(s31[mod*i+2]) , pack(s31[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S32i3 = min_max(pack(s31[mod*i+3]) , pack(s31[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S32i4 = min_max(pack(s31[mod*i+4]) , pack(s31[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S32i5 = min_max(pack(s31[mod*i+5]) , pack(s31[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S32i6 = min_max(pack(s31[mod*i+6]) , pack(s31[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S32i7 = min_max(pack(s31[mod*i+7]) , pack(s31[mod*i+7+mod/2]));
			 Vector#(2, Int#(32)) _S32i8 = min_max(pack(s31[mod*i+8]) , pack(s31[mod*i+8+mod/2]));
			 Vector#(2, Int#(32)) _S32i9 = min_max(pack(s31[mod*i+9]) , pack(s31[mod*i+9+mod/2]));
			 Vector#(2, Int#(32)) _S32i10 = min_max(pack(s31[mod*i+10]) , pack(s31[mod*i+10+mod/2]));
			 Vector#(2, Int#(32)) _S32i11 = min_max(pack(s31[mod*i+11]) , pack(s31[mod*i+11+mod/2]));
			 Vector#(2, Int#(32)) _S32i12 = min_max(pack(s31[mod*i+12]) , pack(s31[mod*i+12+mod/2]));
			 Vector#(2, Int#(32)) _S32i13 = min_max(pack(s31[mod*i+13]) , pack(s31[mod*i+13+mod/2]));
			 Vector#(2, Int#(32)) _S32i14 = min_max(pack(s31[mod*i+14]) , pack(s31[mod*i+14+mod/2]));
			 Vector#(2, Int#(32)) _S32i15 = min_max(pack(s31[mod*i+15]) , pack(s31[mod*i+15+mod/2]));
		if ((i/8)%2 == 0) begin
			s32[mod*i+0] <= _S32i0[0];
			s32[mod*i+0+mod/2] <= _S32i0[1];
			s32[mod*i+1] <= _S32i1[0];
			s32[mod*i+1+mod/2] <= _S32i1[1];
			s32[mod*i+2] <= _S32i2[0];
			s32[mod*i+2+mod/2] <= _S32i2[1];
			s32[mod*i+3] <= _S32i3[0];
			s32[mod*i+3+mod/2] <= _S32i3[1];
			s32[mod*i+4] <= _S32i4[0];
			s32[mod*i+4+mod/2] <= _S32i4[1];
			s32[mod*i+5] <= _S32i5[0];
			s32[mod*i+5+mod/2] <= _S32i5[1];
			s32[mod*i+6] <= _S32i6[0];
			s32[mod*i+6+mod/2] <= _S32i6[1];
			s32[mod*i+7] <= _S32i7[0];
			s32[mod*i+7+mod/2] <= _S32i7[1];
			s32[mod*i+8] <= _S32i8[0];
			s32[mod*i+8+mod/2] <= _S32i8[1];
			s32[mod*i+9] <= _S32i9[0];
			s32[mod*i+9+mod/2] <= _S32i9[1];
			s32[mod*i+10] <= _S32i10[0];
			s32[mod*i+10+mod/2] <= _S32i10[1];
			s32[mod*i+11] <= _S32i11[0];
			s32[mod*i+11+mod/2] <= _S32i11[1];
			s32[mod*i+12] <= _S32i12[0];
			s32[mod*i+12+mod/2] <= _S32i12[1];
			s32[mod*i+13] <= _S32i13[0];
			s32[mod*i+13+mod/2] <= _S32i13[1];
			s32[mod*i+14] <= _S32i14[0];
			s32[mod*i+14+mod/2] <= _S32i14[1];
			s32[mod*i+15] <= _S32i15[0];
			s32[mod*i+15+mod/2] <= _S32i15[1];
		end
		else begin
			s32[mod*i+0] <= _S32i0[1];
			s32[mod*i+0+mod/2] <= _S32i0[0];
			s32[mod*i+1] <= _S32i1[1];
			s32[mod*i+1+mod/2] <= _S32i1[0];
			s32[mod*i+2] <= _S32i2[1];
			s32[mod*i+2+mod/2] <= _S32i2[0];
			s32[mod*i+3] <= _S32i3[1];
			s32[mod*i+3+mod/2] <= _S32i3[0];
			s32[mod*i+4] <= _S32i4[1];
			s32[mod*i+4+mod/2] <= _S32i4[0];
			s32[mod*i+5] <= _S32i5[1];
			s32[mod*i+5+mod/2] <= _S32i5[0];
			s32[mod*i+6] <= _S32i6[1];
			s32[mod*i+6+mod/2] <= _S32i6[0];
			s32[mod*i+7] <= _S32i7[1];
			s32[mod*i+7+mod/2] <= _S32i7[0];
			s32[mod*i+8] <= _S32i8[1];
			s32[mod*i+8+mod/2] <= _S32i8[0];
			s32[mod*i+9] <= _S32i9[1];
			s32[mod*i+9+mod/2] <= _S32i9[0];
			s32[mod*i+10] <= _S32i10[1];
			s32[mod*i+10+mod/2] <= _S32i10[0];
			s32[mod*i+11] <= _S32i11[1];
			s32[mod*i+11+mod/2] <= _S32i11[0];
			s32[mod*i+12] <= _S32i12[1];
			s32[mod*i+12+mod/2] <= _S32i12[0];
			s32[mod*i+13] <= _S32i13[1];
			s32[mod*i+13+mod/2] <= _S32i13[0];
			s32[mod*i+14] <= _S32i14[1];
			s32[mod*i+14+mod/2] <= _S32i14[0];
			s32[mod*i+15] <= _S32i15[1];
			s32[mod*i+15+mod/2] <= _S32i15[0];
		end
	end
	p32.enq(1);
endrule
rule _Q74;
	p32.deq;
	let mod = 16;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S33i0 = min_max(pack(s32[mod*i+0]) , pack(s32[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S33i1 = min_max(pack(s32[mod*i+1]) , pack(s32[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S33i2 = min_max(pack(s32[mod*i+2]) , pack(s32[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S33i3 = min_max(pack(s32[mod*i+3]) , pack(s32[mod*i+3+mod/2]));
			 Vector#(2, Int#(32)) _S33i4 = min_max(pack(s32[mod*i+4]) , pack(s32[mod*i+4+mod/2]));
			 Vector#(2, Int#(32)) _S33i5 = min_max(pack(s32[mod*i+5]) , pack(s32[mod*i+5+mod/2]));
			 Vector#(2, Int#(32)) _S33i6 = min_max(pack(s32[mod*i+6]) , pack(s32[mod*i+6+mod/2]));
			 Vector#(2, Int#(32)) _S33i7 = min_max(pack(s32[mod*i+7]) , pack(s32[mod*i+7+mod/2]));
		if ((i/16)%2 == 0) begin
			s33[mod*i+0] <= _S33i0[0];
			s33[mod*i+0+mod/2] <= _S33i0[1];
			s33[mod*i+1] <= _S33i1[0];
			s33[mod*i+1+mod/2] <= _S33i1[1];
			s33[mod*i+2] <= _S33i2[0];
			s33[mod*i+2+mod/2] <= _S33i2[1];
			s33[mod*i+3] <= _S33i3[0];
			s33[mod*i+3+mod/2] <= _S33i3[1];
			s33[mod*i+4] <= _S33i4[0];
			s33[mod*i+4+mod/2] <= _S33i4[1];
			s33[mod*i+5] <= _S33i5[0];
			s33[mod*i+5+mod/2] <= _S33i5[1];
			s33[mod*i+6] <= _S33i6[0];
			s33[mod*i+6+mod/2] <= _S33i6[1];
			s33[mod*i+7] <= _S33i7[0];
			s33[mod*i+7+mod/2] <= _S33i7[1];
		end
		else begin
			s33[mod*i+0] <= _S33i0[1];
			s33[mod*i+0+mod/2] <= _S33i0[0];
			s33[mod*i+1] <= _S33i1[1];
			s33[mod*i+1+mod/2] <= _S33i1[0];
			s33[mod*i+2] <= _S33i2[1];
			s33[mod*i+2+mod/2] <= _S33i2[0];
			s33[mod*i+3] <= _S33i3[1];
			s33[mod*i+3+mod/2] <= _S33i3[0];
			s33[mod*i+4] <= _S33i4[1];
			s33[mod*i+4+mod/2] <= _S33i4[0];
			s33[mod*i+5] <= _S33i5[1];
			s33[mod*i+5+mod/2] <= _S33i5[0];
			s33[mod*i+6] <= _S33i6[1];
			s33[mod*i+6+mod/2] <= _S33i6[0];
			s33[mod*i+7] <= _S33i7[1];
			s33[mod*i+7+mod/2] <= _S33i7[0];
		end
	end
	p33.enq(1);
endrule
rule _Q73;
	p33.deq;
	let mod = 8;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S34i0 = min_max(pack(s33[mod*i+0]) , pack(s33[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S34i1 = min_max(pack(s33[mod*i+1]) , pack(s33[mod*i+1+mod/2]));
			 Vector#(2, Int#(32)) _S34i2 = min_max(pack(s33[mod*i+2]) , pack(s33[mod*i+2+mod/2]));
			 Vector#(2, Int#(32)) _S34i3 = min_max(pack(s33[mod*i+3]) , pack(s33[mod*i+3+mod/2]));
		if ((i/32)%2 == 0) begin
			s34[mod*i+0] <= _S34i0[0];
			s34[mod*i+0+mod/2] <= _S34i0[1];
			s34[mod*i+1] <= _S34i1[0];
			s34[mod*i+1+mod/2] <= _S34i1[1];
			s34[mod*i+2] <= _S34i2[0];
			s34[mod*i+2+mod/2] <= _S34i2[1];
			s34[mod*i+3] <= _S34i3[0];
			s34[mod*i+3+mod/2] <= _S34i3[1];
		end
		else begin
			s34[mod*i+0] <= _S34i0[1];
			s34[mod*i+0+mod/2] <= _S34i0[0];
			s34[mod*i+1] <= _S34i1[1];
			s34[mod*i+1+mod/2] <= _S34i1[0];
			s34[mod*i+2] <= _S34i2[1];
			s34[mod*i+2+mod/2] <= _S34i2[0];
			s34[mod*i+3] <= _S34i3[1];
			s34[mod*i+3+mod/2] <= _S34i3[0];
		end
	end
	p34.enq(1);
endrule
rule _Q72;
	p34.deq;
	let mod = 4;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S35i0 = min_max(pack(s34[mod*i+0]) , pack(s34[mod*i+0+mod/2]));
			 Vector#(2, Int#(32)) _S35i1 = min_max(pack(s34[mod*i+1]) , pack(s34[mod*i+1+mod/2]));
		if ((i/64)%2 == 0) begin
			s35[mod*i+0] <= _S35i0[0];
			s35[mod*i+0+mod/2] <= _S35i0[1];
			s35[mod*i+1] <= _S35i1[0];
			s35[mod*i+1+mod/2] <= _S35i1[1];
		end
		else begin
			s35[mod*i+0] <= _S35i0[1];
			s35[mod*i+0+mod/2] <= _S35i0[0];
			s35[mod*i+1] <= _S35i1[1];
			s35[mod*i+1+mod/2] <= _S35i1[0];
		end
	end
	p35.enq(1);
endrule
rule _Q71;
	p35.deq;
	let mod = 2;
	for(int i=0; i < L0/mod; i = i + 1) begin
			 Vector#(2, Int#(32)) _S36i0 = min_max(pack(s35[mod*i+0]) , pack(s35[mod*i+0+mod/2]));
		if ((i/128)%2 == 0) begin
			s36[mod*i+0] <= _S36i0[0];
			s36[mod*i+0+mod/2] <= _S36i0[1];
		end
		else begin
			s36[mod*i+0] <= _S36i0[1];
			s36[mod*i+0+mod/2] <= _S36i0[0];
		end
	end
	p36.enq(1);
endrule

method Action put(Vector#(L0, Int#(32)) datas);
for(int i=0;i<L0;i=i+1)
s0[i] <= datas[i];
p0.enq(1);
endmethod

method ActionValue#(Vector#(L0, Int#(32))) get;
p36.deq;
Vector#(L0,Int#(32)) r = newVector;
for(int i=0; i<L0; i = i + 1)
r[i] = s36[i];
return r;
endmethod
endmodule
endpackage