package flowtest;
import FIFO::*;
import FIFOF::*;
import datatypes::*;
import SpecialFIFOs:: * ;
import Real::*;
import Vector::*;
import bitonic::*;
#define L0 128
(*synthesize*)
module mkFlowTest();

Bitonic px <- mkBitonic;

	rule push_data;
		Vector#(L0,Int#(16)) r = newVector;
		for (Int  # (16) i=0; i<L0; i = i + 1)
		r[0]=601;
		r[1]=164;
		r[2]=708;
		r[3]=377;
		r[4]=589;
		r[5]=360;
		r[6]=706;
		r[7]=303;
		r[8]=138;
		r[9]=409;
		r[10]=707;
		r[11]=560;
		r[12]=114;
		r[13]=68;
		r[14]=526;
		r[15]=695;
		r[16]=414;
		r[17]=55;
		r[18]=490;
		r[19]=47;
		r[20]=646;
		r[21]=471;
		r[22]=558;
		r[23]=252;
		r[24]=435;
		r[25]=816;
		r[26]=249;
		r[27]=942;
		r[28]=959;
		r[29]=134;
		r[30]=277;
		r[31]=761;
		r[32]=52;
		r[33]=776;
		r[34]=98;
		r[35]=322;
		r[36]=847;
		r[37]=654;
		r[38]=686;
		r[39]=723;
		r[40]=216;
		r[41]=537;
		r[42]=932;
		r[43]=150;
		r[44]=12;
		r[45]=982;
		r[46]=401;
		r[47]=175;
		r[48]=856;
		r[49]=273;
		r[50]=94;
		r[51]=653;
		r[52]=721;
		r[53]=327;
		r[54]=444;
		r[55]=998;
		r[56]=202;
		r[57]=230;
		r[58]=373;
		r[59]=452;
		r[60]=183;
		r[61]=84;
		r[62]=172;
		r[63]=480;
		r[64]=83;
		r[65]=491;
		r[66]=25;
		r[67]=727;
		r[68]=242;
		r[69]=931;
		r[70]=137;
		r[71]=639;
		r[72]=576;
		r[73]=383;
		r[74]=182;
		r[75]=917;
		r[76]=500;
		r[77]=850;
		r[78]=525;
		r[79]=455;
		r[80]=146;
		r[81]=796;
		r[82]=265;
		r[83]=708;
		r[84]=918;
		r[85]=127;
		r[86]=479;
		r[87]=618;
		r[88]=824;
		r[89]=311;
		r[90]=130;
		r[91]=689;
		r[92]=171;
		r[93]=345;
		r[94]=444;
		r[95]=235;
		r[96]=723;
		r[97]=409;
		r[98]=434;
		r[99]=408;
		r[100]=467;
		r[101]=108;
		r[102]=639;
		r[103]=377;
		r[104]=1000;
		r[105]=772;
		r[106]=898;
		r[107]=865;
		r[108]=362;
		r[109]=62;
		r[110]=346;
		r[111]=204;
		r[112]=712;
		r[113]=80;
		r[114]=37;
		r[115]=275;
		r[116]=807;
		r[117]=142;
		r[118]=941;
		r[119]=740;
		r[120]=386;
		r[121]=281;
		r[122]=959;
		r[123]=693;
		r[124]=975;
		r[125]=149;
		r[126]=350;
		r[127]=518;
		px.put(r);
	endrule


	rule get_data;
	let d <- px.get;
		for(int i=0; i<L0; i=i+1)
			$display("%d",d[i]);
			$finish(0);
	endrule

endmodule
endpackage