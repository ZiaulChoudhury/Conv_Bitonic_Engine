package flowVerilog;
import FixedPoint:: *;
import SpecialFIFOs:: * ;
import Vector:: *;
import FIFO:: *;
import FIFOF:: *;
import datatypes::*;
import compact::*;
#define L0 4096
#define MEMWORD 65536
interface STDIN;
        method Action put(DataType datas);
        method Bit#(16) get;
endinterface

(*synthesize*)
module mkFlowTest(STDIN);
        CompactTree px              <- mkCompactTree;
        Reg#(Int#(16))  cache[L0];
        Reg#(UInt#(12)) sum_count <- mkReg(0);
        Reg#(Int#(16)) total_sum <- mkReg(0);
        Reg#(UInt#(12)) ent <- mkReg(0);
        Reg#(Bit#(MEMWORD)) inQ <- mkReg(0);

        for(int i=0; i < L0; i = i + 1)
                cache[i] <- mkReg(0);
        rule collect (ent == L0);
              px.put(unpack(inQ));
		ent <= 0;
       endrule

        rule receive (sum_count==0);
                let d <- px.get;
		  Vector#(L0,Int#(16)) dx = unpack(d);
                for(int i=0; i < L0; i = i + 1)
                        cache[i] <= dx[i];
                sum_count <= 1;
        endrule
rule s1(sum_count == 1);
  total_sum <= total_sum + cache[0];
endrule
rule s2(sum_count == 2);
  total_sum <= total_sum + cache[1];
endrule
rule s3(sum_count == 3);
  total_sum <= total_sum + cache[2];
endrule
rule s4(sum_count == 4);
  total_sum <= total_sum + cache[3];
endrule
rule s5(sum_count == 5);
  total_sum <= total_sum + cache[4];
endrule
rule s6(sum_count == 6);
  total_sum <= total_sum + cache[5];
endrule
rule s7(sum_count == 7);
  total_sum <= total_sum + cache[6];
endrule
rule s8(sum_count == 8);
  total_sum <= total_sum + cache[7];
endrule
rule s9(sum_count == 9);
  total_sum <= total_sum + cache[8];
endrule
rule s10(sum_count == 10);
  total_sum <= total_sum + cache[9];
endrule
rule s11(sum_count == 11);
  total_sum <= total_sum + cache[10];
endrule
rule s12(sum_count == 12);
  total_sum <= total_sum + cache[11];
endrule
rule s13(sum_count == 13);
  total_sum <= total_sum + cache[12];
endrule
rule s14(sum_count == 14);
  total_sum <= total_sum + cache[13];
endrule
rule s15(sum_count == 15);
  total_sum <= total_sum + cache[14];
endrule
rule s16(sum_count == 16);
  total_sum <= total_sum + cache[15];
endrule
rule s17(sum_count == 17);
  total_sum <= total_sum + cache[16];
endrule
rule s18(sum_count == 18);
  total_sum <= total_sum + cache[17];
endrule
rule s19(sum_count == 19);
  total_sum <= total_sum + cache[18];
endrule
rule s20(sum_count == 20);
  total_sum <= total_sum + cache[19];
endrule
rule s21(sum_count == 21);
  total_sum <= total_sum + cache[20];
endrule
rule s22(sum_count == 22);
  total_sum <= total_sum + cache[21];
endrule
rule s23(sum_count == 23);
  total_sum <= total_sum + cache[22];
endrule
rule s24(sum_count == 24);
  total_sum <= total_sum + cache[23];
endrule
rule s25(sum_count == 25);
  total_sum <= total_sum + cache[24];
endrule
rule s26(sum_count == 26);
  total_sum <= total_sum + cache[25];
endrule
rule s27(sum_count == 27);
  total_sum <= total_sum + cache[26];
endrule
rule s28(sum_count == 28);
  total_sum <= total_sum + cache[27];
endrule
rule s29(sum_count == 29);
  total_sum <= total_sum + cache[28];
endrule
rule s30(sum_count == 30);
  total_sum <= total_sum + cache[29];
endrule
rule s31(sum_count == 31);
  total_sum <= total_sum + cache[30];
endrule
rule s32(sum_count == 32);
  total_sum <= total_sum + cache[31];
endrule
rule s33(sum_count == 33);
  total_sum <= total_sum + cache[32];
endrule
rule s34(sum_count == 34);
  total_sum <= total_sum + cache[33];
endrule
rule s35(sum_count == 35);
  total_sum <= total_sum + cache[34];
endrule
rule s36(sum_count == 36);
  total_sum <= total_sum + cache[35];
endrule
rule s37(sum_count == 37);
  total_sum <= total_sum + cache[36];
endrule
rule s38(sum_count == 38);
  total_sum <= total_sum + cache[37];
endrule
rule s39(sum_count == 39);
  total_sum <= total_sum + cache[38];
endrule
rule s40(sum_count == 40);
  total_sum <= total_sum + cache[39];
endrule
rule s41(sum_count == 41);
  total_sum <= total_sum + cache[40];
endrule
rule s42(sum_count == 42);
  total_sum <= total_sum + cache[41];
endrule
rule s43(sum_count == 43);
  total_sum <= total_sum + cache[42];
endrule
rule s44(sum_count == 44);
  total_sum <= total_sum + cache[43];
endrule
rule s45(sum_count == 45);
  total_sum <= total_sum + cache[44];
endrule
rule s46(sum_count == 46);
  total_sum <= total_sum + cache[45];
endrule
rule s47(sum_count == 47);
  total_sum <= total_sum + cache[46];
endrule
rule s48(sum_count == 48);
  total_sum <= total_sum + cache[47];
endrule
rule s49(sum_count == 49);
  total_sum <= total_sum + cache[48];
endrule
rule s50(sum_count == 50);
  total_sum <= total_sum + cache[49];
endrule
rule s51(sum_count == 51);
  total_sum <= total_sum + cache[50];
endrule
rule s52(sum_count == 52);
  total_sum <= total_sum + cache[51];
endrule
rule s53(sum_count == 53);
  total_sum <= total_sum + cache[52];
endrule
rule s54(sum_count == 54);
  total_sum <= total_sum + cache[53];
endrule
rule s55(sum_count == 55);
  total_sum <= total_sum + cache[54];
endrule
rule s56(sum_count == 56);
  total_sum <= total_sum + cache[55];
endrule
rule s57(sum_count == 57);
  total_sum <= total_sum + cache[56];
endrule
rule s58(sum_count == 58);
  total_sum <= total_sum + cache[57];
endrule
rule s59(sum_count == 59);
  total_sum <= total_sum + cache[58];
endrule
rule s60(sum_count == 60);
  total_sum <= total_sum + cache[59];
endrule
rule s61(sum_count == 61);
  total_sum <= total_sum + cache[60];
endrule
rule s62(sum_count == 62);
  total_sum <= total_sum + cache[61];
endrule
rule s63(sum_count == 63);
  total_sum <= total_sum + cache[62];
endrule
rule s64(sum_count == 64);
  total_sum <= total_sum + cache[63];
endrule
rule s65(sum_count == 65);
  total_sum <= total_sum + cache[64];
endrule
rule s66(sum_count == 66);
  total_sum <= total_sum + cache[65];
endrule
rule s67(sum_count == 67);
  total_sum <= total_sum + cache[66];
endrule
rule s68(sum_count == 68);
  total_sum <= total_sum + cache[67];
endrule
rule s69(sum_count == 69);
  total_sum <= total_sum + cache[68];
endrule
rule s70(sum_count == 70);
  total_sum <= total_sum + cache[69];
endrule
rule s71(sum_count == 71);
  total_sum <= total_sum + cache[70];
endrule
rule s72(sum_count == 72);
  total_sum <= total_sum + cache[71];
endrule
rule s73(sum_count == 73);
  total_sum <= total_sum + cache[72];
endrule
rule s74(sum_count == 74);
  total_sum <= total_sum + cache[73];
endrule
rule s75(sum_count == 75);
  total_sum <= total_sum + cache[74];
endrule
rule s76(sum_count == 76);
  total_sum <= total_sum + cache[75];
endrule
rule s77(sum_count == 77);
  total_sum <= total_sum + cache[76];
endrule
rule s78(sum_count == 78);
  total_sum <= total_sum + cache[77];
endrule
rule s79(sum_count == 79);
  total_sum <= total_sum + cache[78];
endrule
rule s80(sum_count == 80);
  total_sum <= total_sum + cache[79];
endrule
rule s81(sum_count == 81);
  total_sum <= total_sum + cache[80];
endrule
rule s82(sum_count == 82);
  total_sum <= total_sum + cache[81];
endrule
rule s83(sum_count == 83);
  total_sum <= total_sum + cache[82];
endrule
rule s84(sum_count == 84);
  total_sum <= total_sum + cache[83];
endrule
rule s85(sum_count == 85);
  total_sum <= total_sum + cache[84];
endrule
rule s86(sum_count == 86);
  total_sum <= total_sum + cache[85];
endrule
rule s87(sum_count == 87);
  total_sum <= total_sum + cache[86];
endrule
rule s88(sum_count == 88);
  total_sum <= total_sum + cache[87];
endrule
rule s89(sum_count == 89);
  total_sum <= total_sum + cache[88];
endrule
rule s90(sum_count == 90);
  total_sum <= total_sum + cache[89];
endrule
rule s91(sum_count == 91);
  total_sum <= total_sum + cache[90];
endrule
rule s92(sum_count == 92);
  total_sum <= total_sum + cache[91];
endrule
rule s93(sum_count == 93);
  total_sum <= total_sum + cache[92];
endrule
rule s94(sum_count == 94);
  total_sum <= total_sum + cache[93];
endrule
rule s95(sum_count == 95);
  total_sum <= total_sum + cache[94];
endrule
rule s96(sum_count == 96);
  total_sum <= total_sum + cache[95];
endrule
rule s97(sum_count == 97);
  total_sum <= total_sum + cache[96];
endrule
rule s98(sum_count == 98);
  total_sum <= total_sum + cache[97];
endrule
rule s99(sum_count == 99);
  total_sum <= total_sum + cache[98];
endrule
rule s100(sum_count == 100);
  total_sum <= total_sum + cache[99];
endrule
rule s101(sum_count == 101);
  total_sum <= total_sum + cache[100];
endrule
rule s102(sum_count == 102);
  total_sum <= total_sum + cache[101];
endrule
rule s103(sum_count == 103);
  total_sum <= total_sum + cache[102];
endrule
rule s104(sum_count == 104);
  total_sum <= total_sum + cache[103];
endrule
rule s105(sum_count == 105);
  total_sum <= total_sum + cache[104];
endrule
rule s106(sum_count == 106);
  total_sum <= total_sum + cache[105];
endrule
rule s107(sum_count == 107);
  total_sum <= total_sum + cache[106];
endrule
rule s108(sum_count == 108);
  total_sum <= total_sum + cache[107];
endrule
rule s109(sum_count == 109);
  total_sum <= total_sum + cache[108];
endrule
rule s110(sum_count == 110);
  total_sum <= total_sum + cache[109];
endrule
rule s111(sum_count == 111);
  total_sum <= total_sum + cache[110];
endrule
rule s112(sum_count == 112);
  total_sum <= total_sum + cache[111];
endrule
rule s113(sum_count == 113);
  total_sum <= total_sum + cache[112];
endrule
rule s114(sum_count == 114);
  total_sum <= total_sum + cache[113];
endrule
rule s115(sum_count == 115);
  total_sum <= total_sum + cache[114];
endrule
rule s116(sum_count == 116);
  total_sum <= total_sum + cache[115];
endrule
rule s117(sum_count == 117);
  total_sum <= total_sum + cache[116];
endrule
rule s118(sum_count == 118);
  total_sum <= total_sum + cache[117];
endrule
rule s119(sum_count == 119);
  total_sum <= total_sum + cache[118];
endrule
rule s120(sum_count == 120);
  total_sum <= total_sum + cache[119];
endrule
rule s121(sum_count == 121);
  total_sum <= total_sum + cache[120];
endrule
rule s122(sum_count == 122);
  total_sum <= total_sum + cache[121];
endrule
rule s123(sum_count == 123);
  total_sum <= total_sum + cache[122];
endrule
rule s124(sum_count == 124);
  total_sum <= total_sum + cache[123];
endrule
rule s125(sum_count == 125);
  total_sum <= total_sum + cache[124];
endrule
rule s126(sum_count == 126);
  total_sum <= total_sum + cache[125];
endrule
rule s127(sum_count == 127);
  total_sum <= total_sum + cache[126];
endrule
rule s128(sum_count == 128);
  total_sum <= total_sum + cache[127];
endrule
rule s129(sum_count == 129);
  total_sum <= total_sum + cache[128];
endrule
rule s130(sum_count == 130);
  total_sum <= total_sum + cache[129];
endrule
rule s131(sum_count == 131);
  total_sum <= total_sum + cache[130];
endrule
rule s132(sum_count == 132);
  total_sum <= total_sum + cache[131];
endrule
rule s133(sum_count == 133);
  total_sum <= total_sum + cache[132];
endrule
rule s134(sum_count == 134);
  total_sum <= total_sum + cache[133];
endrule
rule s135(sum_count == 135);
  total_sum <= total_sum + cache[134];
endrule
rule s136(sum_count == 136);
  total_sum <= total_sum + cache[135];
endrule
rule s137(sum_count == 137);
  total_sum <= total_sum + cache[136];
endrule
rule s138(sum_count == 138);
  total_sum <= total_sum + cache[137];
endrule
rule s139(sum_count == 139);
  total_sum <= total_sum + cache[138];
endrule
rule s140(sum_count == 140);
  total_sum <= total_sum + cache[139];
endrule
rule s141(sum_count == 141);
  total_sum <= total_sum + cache[140];
endrule
rule s142(sum_count == 142);
  total_sum <= total_sum + cache[141];
endrule
rule s143(sum_count == 143);
  total_sum <= total_sum + cache[142];
endrule
rule s144(sum_count == 144);
  total_sum <= total_sum + cache[143];
endrule
rule s145(sum_count == 145);
  total_sum <= total_sum + cache[144];
endrule
rule s146(sum_count == 146);
  total_sum <= total_sum + cache[145];
endrule
rule s147(sum_count == 147);
  total_sum <= total_sum + cache[146];
endrule
rule s148(sum_count == 148);
  total_sum <= total_sum + cache[147];
endrule
rule s149(sum_count == 149);
  total_sum <= total_sum + cache[148];
endrule
rule s150(sum_count == 150);
  total_sum <= total_sum + cache[149];
endrule
rule s151(sum_count == 151);
  total_sum <= total_sum + cache[150];
endrule
rule s152(sum_count == 152);
  total_sum <= total_sum + cache[151];
endrule
rule s153(sum_count == 153);
  total_sum <= total_sum + cache[152];
endrule
rule s154(sum_count == 154);
  total_sum <= total_sum + cache[153];
endrule
rule s155(sum_count == 155);
  total_sum <= total_sum + cache[154];
endrule
rule s156(sum_count == 156);
  total_sum <= total_sum + cache[155];
endrule
rule s157(sum_count == 157);
  total_sum <= total_sum + cache[156];
endrule
rule s158(sum_count == 158);
  total_sum <= total_sum + cache[157];
endrule
rule s159(sum_count == 159);
  total_sum <= total_sum + cache[158];
endrule
rule s160(sum_count == 160);
  total_sum <= total_sum + cache[159];
endrule
rule s161(sum_count == 161);
  total_sum <= total_sum + cache[160];
endrule
rule s162(sum_count == 162);
  total_sum <= total_sum + cache[161];
endrule
rule s163(sum_count == 163);
  total_sum <= total_sum + cache[162];
endrule
rule s164(sum_count == 164);
  total_sum <= total_sum + cache[163];
endrule
rule s165(sum_count == 165);
  total_sum <= total_sum + cache[164];
endrule
rule s166(sum_count == 166);
  total_sum <= total_sum + cache[165];
endrule
rule s167(sum_count == 167);
  total_sum <= total_sum + cache[166];
endrule
rule s168(sum_count == 168);
  total_sum <= total_sum + cache[167];
endrule
rule s169(sum_count == 169);
  total_sum <= total_sum + cache[168];
endrule
rule s170(sum_count == 170);
  total_sum <= total_sum + cache[169];
endrule
rule s171(sum_count == 171);
  total_sum <= total_sum + cache[170];
endrule
rule s172(sum_count == 172);
  total_sum <= total_sum + cache[171];
endrule
rule s173(sum_count == 173);
  total_sum <= total_sum + cache[172];
endrule
rule s174(sum_count == 174);
  total_sum <= total_sum + cache[173];
endrule
rule s175(sum_count == 175);
  total_sum <= total_sum + cache[174];
endrule
rule s176(sum_count == 176);
  total_sum <= total_sum + cache[175];
endrule
rule s177(sum_count == 177);
  total_sum <= total_sum + cache[176];
endrule
rule s178(sum_count == 178);
  total_sum <= total_sum + cache[177];
endrule
rule s179(sum_count == 179);
  total_sum <= total_sum + cache[178];
endrule
rule s180(sum_count == 180);
  total_sum <= total_sum + cache[179];
endrule
rule s181(sum_count == 181);
  total_sum <= total_sum + cache[180];
endrule
rule s182(sum_count == 182);
  total_sum <= total_sum + cache[181];
endrule
rule s183(sum_count == 183);
  total_sum <= total_sum + cache[182];
endrule
rule s184(sum_count == 184);
  total_sum <= total_sum + cache[183];
endrule
rule s185(sum_count == 185);
  total_sum <= total_sum + cache[184];
endrule
rule s186(sum_count == 186);
  total_sum <= total_sum + cache[185];
endrule
rule s187(sum_count == 187);
  total_sum <= total_sum + cache[186];
endrule
rule s188(sum_count == 188);
  total_sum <= total_sum + cache[187];
endrule
rule s189(sum_count == 189);
  total_sum <= total_sum + cache[188];
endrule
rule s190(sum_count == 190);
  total_sum <= total_sum + cache[189];
endrule
rule s191(sum_count == 191);
  total_sum <= total_sum + cache[190];
endrule
rule s192(sum_count == 192);
  total_sum <= total_sum + cache[191];
endrule
rule s193(sum_count == 193);
  total_sum <= total_sum + cache[192];
endrule
rule s194(sum_count == 194);
  total_sum <= total_sum + cache[193];
endrule
rule s195(sum_count == 195);
  total_sum <= total_sum + cache[194];
endrule
rule s196(sum_count == 196);
  total_sum <= total_sum + cache[195];
endrule
rule s197(sum_count == 197);
  total_sum <= total_sum + cache[196];
endrule
rule s198(sum_count == 198);
  total_sum <= total_sum + cache[197];
endrule
rule s199(sum_count == 199);
  total_sum <= total_sum + cache[198];
endrule
rule s200(sum_count == 200);
  total_sum <= total_sum + cache[199];
endrule
rule s201(sum_count == 201);
  total_sum <= total_sum + cache[200];
endrule
rule s202(sum_count == 202);
  total_sum <= total_sum + cache[201];
endrule
rule s203(sum_count == 203);
  total_sum <= total_sum + cache[202];
endrule
rule s204(sum_count == 204);
  total_sum <= total_sum + cache[203];
endrule
rule s205(sum_count == 205);
  total_sum <= total_sum + cache[204];
endrule
rule s206(sum_count == 206);
  total_sum <= total_sum + cache[205];
endrule
rule s207(sum_count == 207);
  total_sum <= total_sum + cache[206];
endrule
rule s208(sum_count == 208);
  total_sum <= total_sum + cache[207];
endrule
rule s209(sum_count == 209);
  total_sum <= total_sum + cache[208];
endrule
rule s210(sum_count == 210);
  total_sum <= total_sum + cache[209];
endrule
rule s211(sum_count == 211);
  total_sum <= total_sum + cache[210];
endrule
rule s212(sum_count == 212);
  total_sum <= total_sum + cache[211];
endrule
rule s213(sum_count == 213);
  total_sum <= total_sum + cache[212];
endrule
rule s214(sum_count == 214);
  total_sum <= total_sum + cache[213];
endrule
rule s215(sum_count == 215);
  total_sum <= total_sum + cache[214];
endrule
rule s216(sum_count == 216);
  total_sum <= total_sum + cache[215];
endrule
rule s217(sum_count == 217);
  total_sum <= total_sum + cache[216];
endrule
rule s218(sum_count == 218);
  total_sum <= total_sum + cache[217];
endrule
rule s219(sum_count == 219);
  total_sum <= total_sum + cache[218];
endrule
rule s220(sum_count == 220);
  total_sum <= total_sum + cache[219];
endrule
rule s221(sum_count == 221);
  total_sum <= total_sum + cache[220];
endrule
rule s222(sum_count == 222);
  total_sum <= total_sum + cache[221];
endrule
rule s223(sum_count == 223);
  total_sum <= total_sum + cache[222];
endrule
rule s224(sum_count == 224);
  total_sum <= total_sum + cache[223];
endrule
rule s225(sum_count == 225);
  total_sum <= total_sum + cache[224];
endrule
rule s226(sum_count == 226);
  total_sum <= total_sum + cache[225];
endrule
rule s227(sum_count == 227);
  total_sum <= total_sum + cache[226];
endrule
rule s228(sum_count == 228);
  total_sum <= total_sum + cache[227];
endrule
rule s229(sum_count == 229);
  total_sum <= total_sum + cache[228];
endrule
rule s230(sum_count == 230);
  total_sum <= total_sum + cache[229];
endrule
rule s231(sum_count == 231);
  total_sum <= total_sum + cache[230];
endrule
rule s232(sum_count == 232);
  total_sum <= total_sum + cache[231];
endrule
rule s233(sum_count == 233);
  total_sum <= total_sum + cache[232];
endrule
rule s234(sum_count == 234);
  total_sum <= total_sum + cache[233];
endrule
rule s235(sum_count == 235);
  total_sum <= total_sum + cache[234];
endrule
rule s236(sum_count == 236);
  total_sum <= total_sum + cache[235];
endrule
rule s237(sum_count == 237);
  total_sum <= total_sum + cache[236];
endrule
rule s238(sum_count == 238);
  total_sum <= total_sum + cache[237];
endrule
rule s239(sum_count == 239);
  total_sum <= total_sum + cache[238];
endrule
rule s240(sum_count == 240);
  total_sum <= total_sum + cache[239];
endrule
rule s241(sum_count == 241);
  total_sum <= total_sum + cache[240];
endrule
rule s242(sum_count == 242);
  total_sum <= total_sum + cache[241];
endrule
rule s243(sum_count == 243);
  total_sum <= total_sum + cache[242];
endrule
rule s244(sum_count == 244);
  total_sum <= total_sum + cache[243];
endrule
rule s245(sum_count == 245);
  total_sum <= total_sum + cache[244];
endrule
rule s246(sum_count == 246);
  total_sum <= total_sum + cache[245];
endrule
rule s247(sum_count == 247);
  total_sum <= total_sum + cache[246];
endrule
rule s248(sum_count == 248);
  total_sum <= total_sum + cache[247];
endrule
rule s249(sum_count == 249);
  total_sum <= total_sum + cache[248];
endrule
rule s250(sum_count == 250);
  total_sum <= total_sum + cache[249];
endrule
rule s251(sum_count == 251);
  total_sum <= total_sum + cache[250];
endrule
rule s252(sum_count == 252);
  total_sum <= total_sum + cache[251];
endrule
rule s253(sum_count == 253);
  total_sum <= total_sum + cache[252];
endrule
rule s254(sum_count == 254);
  total_sum <= total_sum + cache[253];
endrule
rule s255(sum_count == 255);
  total_sum <= total_sum + cache[254];
endrule
rule s256(sum_count == 256);
  total_sum <= total_sum + cache[255];
endrule
rule s257(sum_count == 257);
  total_sum <= total_sum + cache[256];
endrule
rule s258(sum_count == 258);
  total_sum <= total_sum + cache[257];
endrule
rule s259(sum_count == 259);
  total_sum <= total_sum + cache[258];
endrule
rule s260(sum_count == 260);
  total_sum <= total_sum + cache[259];
endrule
rule s261(sum_count == 261);
  total_sum <= total_sum + cache[260];
endrule
rule s262(sum_count == 262);
  total_sum <= total_sum + cache[261];
endrule
rule s263(sum_count == 263);
  total_sum <= total_sum + cache[262];
endrule
rule s264(sum_count == 264);
  total_sum <= total_sum + cache[263];
endrule
rule s265(sum_count == 265);
  total_sum <= total_sum + cache[264];
endrule
rule s266(sum_count == 266);
  total_sum <= total_sum + cache[265];
endrule
rule s267(sum_count == 267);
  total_sum <= total_sum + cache[266];
endrule
rule s268(sum_count == 268);
  total_sum <= total_sum + cache[267];
endrule
rule s269(sum_count == 269);
  total_sum <= total_sum + cache[268];
endrule
rule s270(sum_count == 270);
  total_sum <= total_sum + cache[269];
endrule
rule s271(sum_count == 271);
  total_sum <= total_sum + cache[270];
endrule
rule s272(sum_count == 272);
  total_sum <= total_sum + cache[271];
endrule
rule s273(sum_count == 273);
  total_sum <= total_sum + cache[272];
endrule
rule s274(sum_count == 274);
  total_sum <= total_sum + cache[273];
endrule
rule s275(sum_count == 275);
  total_sum <= total_sum + cache[274];
endrule
rule s276(sum_count == 276);
  total_sum <= total_sum + cache[275];
endrule
rule s277(sum_count == 277);
  total_sum <= total_sum + cache[276];
endrule
rule s278(sum_count == 278);
  total_sum <= total_sum + cache[277];
endrule
rule s279(sum_count == 279);
  total_sum <= total_sum + cache[278];
endrule
rule s280(sum_count == 280);
  total_sum <= total_sum + cache[279];
endrule
rule s281(sum_count == 281);
  total_sum <= total_sum + cache[280];
endrule
rule s282(sum_count == 282);
  total_sum <= total_sum + cache[281];
endrule
rule s283(sum_count == 283);
  total_sum <= total_sum + cache[282];
endrule
rule s284(sum_count == 284);
  total_sum <= total_sum + cache[283];
endrule
rule s285(sum_count == 285);
  total_sum <= total_sum + cache[284];
endrule
rule s286(sum_count == 286);
  total_sum <= total_sum + cache[285];
endrule
rule s287(sum_count == 287);
  total_sum <= total_sum + cache[286];
endrule
rule s288(sum_count == 288);
  total_sum <= total_sum + cache[287];
endrule
rule s289(sum_count == 289);
  total_sum <= total_sum + cache[288];
endrule
rule s290(sum_count == 290);
  total_sum <= total_sum + cache[289];
endrule
rule s291(sum_count == 291);
  total_sum <= total_sum + cache[290];
endrule
rule s292(sum_count == 292);
  total_sum <= total_sum + cache[291];
endrule
rule s293(sum_count == 293);
  total_sum <= total_sum + cache[292];
endrule
rule s294(sum_count == 294);
  total_sum <= total_sum + cache[293];
endrule
rule s295(sum_count == 295);
  total_sum <= total_sum + cache[294];
endrule
rule s296(sum_count == 296);
  total_sum <= total_sum + cache[295];
endrule
rule s297(sum_count == 297);
  total_sum <= total_sum + cache[296];
endrule
rule s298(sum_count == 298);
  total_sum <= total_sum + cache[297];
endrule
rule s299(sum_count == 299);
  total_sum <= total_sum + cache[298];
endrule
rule s300(sum_count == 300);
  total_sum <= total_sum + cache[299];
endrule
rule s301(sum_count == 301);
  total_sum <= total_sum + cache[300];
endrule
rule s302(sum_count == 302);
  total_sum <= total_sum + cache[301];
endrule
rule s303(sum_count == 303);
  total_sum <= total_sum + cache[302];
endrule
rule s304(sum_count == 304);
  total_sum <= total_sum + cache[303];
endrule
rule s305(sum_count == 305);
  total_sum <= total_sum + cache[304];
endrule
rule s306(sum_count == 306);
  total_sum <= total_sum + cache[305];
endrule
rule s307(sum_count == 307);
  total_sum <= total_sum + cache[306];
endrule
rule s308(sum_count == 308);
  total_sum <= total_sum + cache[307];
endrule
rule s309(sum_count == 309);
  total_sum <= total_sum + cache[308];
endrule
rule s310(sum_count == 310);
  total_sum <= total_sum + cache[309];
endrule
rule s311(sum_count == 311);
  total_sum <= total_sum + cache[310];
endrule
rule s312(sum_count == 312);
  total_sum <= total_sum + cache[311];
endrule
rule s313(sum_count == 313);
  total_sum <= total_sum + cache[312];
endrule
rule s314(sum_count == 314);
  total_sum <= total_sum + cache[313];
endrule
rule s315(sum_count == 315);
  total_sum <= total_sum + cache[314];
endrule
rule s316(sum_count == 316);
  total_sum <= total_sum + cache[315];
endrule
rule s317(sum_count == 317);
  total_sum <= total_sum + cache[316];
endrule
rule s318(sum_count == 318);
  total_sum <= total_sum + cache[317];
endrule
rule s319(sum_count == 319);
  total_sum <= total_sum + cache[318];
endrule
rule s320(sum_count == 320);
  total_sum <= total_sum + cache[319];
endrule
rule s321(sum_count == 321);
  total_sum <= total_sum + cache[320];
endrule
rule s322(sum_count == 322);
  total_sum <= total_sum + cache[321];
endrule
rule s323(sum_count == 323);
  total_sum <= total_sum + cache[322];
endrule
rule s324(sum_count == 324);
  total_sum <= total_sum + cache[323];
endrule
rule s325(sum_count == 325);
  total_sum <= total_sum + cache[324];
endrule
rule s326(sum_count == 326);
  total_sum <= total_sum + cache[325];
endrule
rule s327(sum_count == 327);
  total_sum <= total_sum + cache[326];
endrule
rule s328(sum_count == 328);
  total_sum <= total_sum + cache[327];
endrule
rule s329(sum_count == 329);
  total_sum <= total_sum + cache[328];
endrule
rule s330(sum_count == 330);
  total_sum <= total_sum + cache[329];
endrule
rule s331(sum_count == 331);
  total_sum <= total_sum + cache[330];
endrule
rule s332(sum_count == 332);
  total_sum <= total_sum + cache[331];
endrule
rule s333(sum_count == 333);
  total_sum <= total_sum + cache[332];
endrule
rule s334(sum_count == 334);
  total_sum <= total_sum + cache[333];
endrule
rule s335(sum_count == 335);
  total_sum <= total_sum + cache[334];
endrule
rule s336(sum_count == 336);
  total_sum <= total_sum + cache[335];
endrule
rule s337(sum_count == 337);
  total_sum <= total_sum + cache[336];
endrule
rule s338(sum_count == 338);
  total_sum <= total_sum + cache[337];
endrule
rule s339(sum_count == 339);
  total_sum <= total_sum + cache[338];
endrule
rule s340(sum_count == 340);
  total_sum <= total_sum + cache[339];
endrule
rule s341(sum_count == 341);
  total_sum <= total_sum + cache[340];
endrule
rule s342(sum_count == 342);
  total_sum <= total_sum + cache[341];
endrule
rule s343(sum_count == 343);
  total_sum <= total_sum + cache[342];
endrule
rule s344(sum_count == 344);
  total_sum <= total_sum + cache[343];
endrule
rule s345(sum_count == 345);
  total_sum <= total_sum + cache[344];
endrule
rule s346(sum_count == 346);
  total_sum <= total_sum + cache[345];
endrule
rule s347(sum_count == 347);
  total_sum <= total_sum + cache[346];
endrule
rule s348(sum_count == 348);
  total_sum <= total_sum + cache[347];
endrule
rule s349(sum_count == 349);
  total_sum <= total_sum + cache[348];
endrule
rule s350(sum_count == 350);
  total_sum <= total_sum + cache[349];
endrule
rule s351(sum_count == 351);
  total_sum <= total_sum + cache[350];
endrule
rule s352(sum_count == 352);
  total_sum <= total_sum + cache[351];
endrule
rule s353(sum_count == 353);
  total_sum <= total_sum + cache[352];
endrule
rule s354(sum_count == 354);
  total_sum <= total_sum + cache[353];
endrule
rule s355(sum_count == 355);
  total_sum <= total_sum + cache[354];
endrule
rule s356(sum_count == 356);
  total_sum <= total_sum + cache[355];
endrule
rule s357(sum_count == 357);
  total_sum <= total_sum + cache[356];
endrule
rule s358(sum_count == 358);
  total_sum <= total_sum + cache[357];
endrule
rule s359(sum_count == 359);
  total_sum <= total_sum + cache[358];
endrule
rule s360(sum_count == 360);
  total_sum <= total_sum + cache[359];
endrule
rule s361(sum_count == 361);
  total_sum <= total_sum + cache[360];
endrule
rule s362(sum_count == 362);
  total_sum <= total_sum + cache[361];
endrule
rule s363(sum_count == 363);
  total_sum <= total_sum + cache[362];
endrule
rule s364(sum_count == 364);
  total_sum <= total_sum + cache[363];
endrule
rule s365(sum_count == 365);
  total_sum <= total_sum + cache[364];
endrule
rule s366(sum_count == 366);
  total_sum <= total_sum + cache[365];
endrule
rule s367(sum_count == 367);
  total_sum <= total_sum + cache[366];
endrule
rule s368(sum_count == 368);
  total_sum <= total_sum + cache[367];
endrule
rule s369(sum_count == 369);
  total_sum <= total_sum + cache[368];
endrule
rule s370(sum_count == 370);
  total_sum <= total_sum + cache[369];
endrule
rule s371(sum_count == 371);
  total_sum <= total_sum + cache[370];
endrule
rule s372(sum_count == 372);
  total_sum <= total_sum + cache[371];
endrule
rule s373(sum_count == 373);
  total_sum <= total_sum + cache[372];
endrule
rule s374(sum_count == 374);
  total_sum <= total_sum + cache[373];
endrule
rule s375(sum_count == 375);
  total_sum <= total_sum + cache[374];
endrule
rule s376(sum_count == 376);
  total_sum <= total_sum + cache[375];
endrule
rule s377(sum_count == 377);
  total_sum <= total_sum + cache[376];
endrule
rule s378(sum_count == 378);
  total_sum <= total_sum + cache[377];
endrule
rule s379(sum_count == 379);
  total_sum <= total_sum + cache[378];
endrule
rule s380(sum_count == 380);
  total_sum <= total_sum + cache[379];
endrule
rule s381(sum_count == 381);
  total_sum <= total_sum + cache[380];
endrule
rule s382(sum_count == 382);
  total_sum <= total_sum + cache[381];
endrule
rule s383(sum_count == 383);
  total_sum <= total_sum + cache[382];
endrule
rule s384(sum_count == 384);
  total_sum <= total_sum + cache[383];
endrule
rule s385(sum_count == 385);
  total_sum <= total_sum + cache[384];
endrule
rule s386(sum_count == 386);
  total_sum <= total_sum + cache[385];
endrule
rule s387(sum_count == 387);
  total_sum <= total_sum + cache[386];
endrule
rule s388(sum_count == 388);
  total_sum <= total_sum + cache[387];
endrule
rule s389(sum_count == 389);
  total_sum <= total_sum + cache[388];
endrule
rule s390(sum_count == 390);
  total_sum <= total_sum + cache[389];
endrule
rule s391(sum_count == 391);
  total_sum <= total_sum + cache[390];
endrule
rule s392(sum_count == 392);
  total_sum <= total_sum + cache[391];
endrule
rule s393(sum_count == 393);
  total_sum <= total_sum + cache[392];
endrule
rule s394(sum_count == 394);
  total_sum <= total_sum + cache[393];
endrule
rule s395(sum_count == 395);
  total_sum <= total_sum + cache[394];
endrule
rule s396(sum_count == 396);
  total_sum <= total_sum + cache[395];
endrule
rule s397(sum_count == 397);
  total_sum <= total_sum + cache[396];
endrule
rule s398(sum_count == 398);
  total_sum <= total_sum + cache[397];
endrule
rule s399(sum_count == 399);
  total_sum <= total_sum + cache[398];
endrule
rule s400(sum_count == 400);
  total_sum <= total_sum + cache[399];
endrule
rule s401(sum_count == 401);
  total_sum <= total_sum + cache[400];
endrule
rule s402(sum_count == 402);
  total_sum <= total_sum + cache[401];
endrule
rule s403(sum_count == 403);
  total_sum <= total_sum + cache[402];
endrule
rule s404(sum_count == 404);
  total_sum <= total_sum + cache[403];
endrule
rule s405(sum_count == 405);
  total_sum <= total_sum + cache[404];
endrule
rule s406(sum_count == 406);
  total_sum <= total_sum + cache[405];
endrule
rule s407(sum_count == 407);
  total_sum <= total_sum + cache[406];
endrule
rule s408(sum_count == 408);
  total_sum <= total_sum + cache[407];
endrule
rule s409(sum_count == 409);
  total_sum <= total_sum + cache[408];
endrule
rule s410(sum_count == 410);
  total_sum <= total_sum + cache[409];
endrule
rule s411(sum_count == 411);
  total_sum <= total_sum + cache[410];
endrule
rule s412(sum_count == 412);
  total_sum <= total_sum + cache[411];
endrule
rule s413(sum_count == 413);
  total_sum <= total_sum + cache[412];
endrule
rule s414(sum_count == 414);
  total_sum <= total_sum + cache[413];
endrule
rule s415(sum_count == 415);
  total_sum <= total_sum + cache[414];
endrule
rule s416(sum_count == 416);
  total_sum <= total_sum + cache[415];
endrule
rule s417(sum_count == 417);
  total_sum <= total_sum + cache[416];
endrule
rule s418(sum_count == 418);
  total_sum <= total_sum + cache[417];
endrule
rule s419(sum_count == 419);
  total_sum <= total_sum + cache[418];
endrule
rule s420(sum_count == 420);
  total_sum <= total_sum + cache[419];
endrule
rule s421(sum_count == 421);
  total_sum <= total_sum + cache[420];
endrule
rule s422(sum_count == 422);
  total_sum <= total_sum + cache[421];
endrule
rule s423(sum_count == 423);
  total_sum <= total_sum + cache[422];
endrule
rule s424(sum_count == 424);
  total_sum <= total_sum + cache[423];
endrule
rule s425(sum_count == 425);
  total_sum <= total_sum + cache[424];
endrule
rule s426(sum_count == 426);
  total_sum <= total_sum + cache[425];
endrule
rule s427(sum_count == 427);
  total_sum <= total_sum + cache[426];
endrule
rule s428(sum_count == 428);
  total_sum <= total_sum + cache[427];
endrule
rule s429(sum_count == 429);
  total_sum <= total_sum + cache[428];
endrule
rule s430(sum_count == 430);
  total_sum <= total_sum + cache[429];
endrule
rule s431(sum_count == 431);
  total_sum <= total_sum + cache[430];
endrule
rule s432(sum_count == 432);
  total_sum <= total_sum + cache[431];
endrule
rule s433(sum_count == 433);
  total_sum <= total_sum + cache[432];
endrule
rule s434(sum_count == 434);
  total_sum <= total_sum + cache[433];
endrule
rule s435(sum_count == 435);
  total_sum <= total_sum + cache[434];
endrule
rule s436(sum_count == 436);
  total_sum <= total_sum + cache[435];
endrule
rule s437(sum_count == 437);
  total_sum <= total_sum + cache[436];
endrule
rule s438(sum_count == 438);
  total_sum <= total_sum + cache[437];
endrule
rule s439(sum_count == 439);
  total_sum <= total_sum + cache[438];
endrule
rule s440(sum_count == 440);
  total_sum <= total_sum + cache[439];
endrule
rule s441(sum_count == 441);
  total_sum <= total_sum + cache[440];
endrule
rule s442(sum_count == 442);
  total_sum <= total_sum + cache[441];
endrule
rule s443(sum_count == 443);
  total_sum <= total_sum + cache[442];
endrule
rule s444(sum_count == 444);
  total_sum <= total_sum + cache[443];
endrule
rule s445(sum_count == 445);
  total_sum <= total_sum + cache[444];
endrule
rule s446(sum_count == 446);
  total_sum <= total_sum + cache[445];
endrule
rule s447(sum_count == 447);
  total_sum <= total_sum + cache[446];
endrule
rule s448(sum_count == 448);
  total_sum <= total_sum + cache[447];
endrule
rule s449(sum_count == 449);
  total_sum <= total_sum + cache[448];
endrule
rule s450(sum_count == 450);
  total_sum <= total_sum + cache[449];
endrule
rule s451(sum_count == 451);
  total_sum <= total_sum + cache[450];
endrule
rule s452(sum_count == 452);
  total_sum <= total_sum + cache[451];
endrule
rule s453(sum_count == 453);
  total_sum <= total_sum + cache[452];
endrule
rule s454(sum_count == 454);
  total_sum <= total_sum + cache[453];
endrule
rule s455(sum_count == 455);
  total_sum <= total_sum + cache[454];
endrule
rule s456(sum_count == 456);
  total_sum <= total_sum + cache[455];
endrule
rule s457(sum_count == 457);
  total_sum <= total_sum + cache[456];
endrule
rule s458(sum_count == 458);
  total_sum <= total_sum + cache[457];
endrule
rule s459(sum_count == 459);
  total_sum <= total_sum + cache[458];
endrule
rule s460(sum_count == 460);
  total_sum <= total_sum + cache[459];
endrule
rule s461(sum_count == 461);
  total_sum <= total_sum + cache[460];
endrule
rule s462(sum_count == 462);
  total_sum <= total_sum + cache[461];
endrule
rule s463(sum_count == 463);
  total_sum <= total_sum + cache[462];
endrule
rule s464(sum_count == 464);
  total_sum <= total_sum + cache[463];
endrule
rule s465(sum_count == 465);
  total_sum <= total_sum + cache[464];
endrule
rule s466(sum_count == 466);
  total_sum <= total_sum + cache[465];
endrule
rule s467(sum_count == 467);
  total_sum <= total_sum + cache[466];
endrule
rule s468(sum_count == 468);
  total_sum <= total_sum + cache[467];
endrule
rule s469(sum_count == 469);
  total_sum <= total_sum + cache[468];
endrule
rule s470(sum_count == 470);
  total_sum <= total_sum + cache[469];
endrule
rule s471(sum_count == 471);
  total_sum <= total_sum + cache[470];
endrule
rule s472(sum_count == 472);
  total_sum <= total_sum + cache[471];
endrule
rule s473(sum_count == 473);
  total_sum <= total_sum + cache[472];
endrule
rule s474(sum_count == 474);
  total_sum <= total_sum + cache[473];
endrule
rule s475(sum_count == 475);
  total_sum <= total_sum + cache[474];
endrule
rule s476(sum_count == 476);
  total_sum <= total_sum + cache[475];
endrule
rule s477(sum_count == 477);
  total_sum <= total_sum + cache[476];
endrule
rule s478(sum_count == 478);
  total_sum <= total_sum + cache[477];
endrule
rule s479(sum_count == 479);
  total_sum <= total_sum + cache[478];
endrule
rule s480(sum_count == 480);
  total_sum <= total_sum + cache[479];
endrule
rule s481(sum_count == 481);
  total_sum <= total_sum + cache[480];
endrule
rule s482(sum_count == 482);
  total_sum <= total_sum + cache[481];
endrule
rule s483(sum_count == 483);
  total_sum <= total_sum + cache[482];
endrule
rule s484(sum_count == 484);
  total_sum <= total_sum + cache[483];
endrule
rule s485(sum_count == 485);
  total_sum <= total_sum + cache[484];
endrule
rule s486(sum_count == 486);
  total_sum <= total_sum + cache[485];
endrule
rule s487(sum_count == 487);
  total_sum <= total_sum + cache[486];
endrule
rule s488(sum_count == 488);
  total_sum <= total_sum + cache[487];
endrule
rule s489(sum_count == 489);
  total_sum <= total_sum + cache[488];
endrule
rule s490(sum_count == 490);
  total_sum <= total_sum + cache[489];
endrule
rule s491(sum_count == 491);
  total_sum <= total_sum + cache[490];
endrule
rule s492(sum_count == 492);
  total_sum <= total_sum + cache[491];
endrule
rule s493(sum_count == 493);
  total_sum <= total_sum + cache[492];
endrule
rule s494(sum_count == 494);
  total_sum <= total_sum + cache[493];
endrule
rule s495(sum_count == 495);
  total_sum <= total_sum + cache[494];
endrule
rule s496(sum_count == 496);
  total_sum <= total_sum + cache[495];
endrule
rule s497(sum_count == 497);
  total_sum <= total_sum + cache[496];
endrule
rule s498(sum_count == 498);
  total_sum <= total_sum + cache[497];
endrule
rule s499(sum_count == 499);
  total_sum <= total_sum + cache[498];
endrule
rule s500(sum_count == 500);
  total_sum <= total_sum + cache[499];
endrule
rule s501(sum_count == 501);
  total_sum <= total_sum + cache[500];
endrule
rule s502(sum_count == 502);
  total_sum <= total_sum + cache[501];
endrule
rule s503(sum_count == 503);
  total_sum <= total_sum + cache[502];
endrule
rule s504(sum_count == 504);
  total_sum <= total_sum + cache[503];
endrule
rule s505(sum_count == 505);
  total_sum <= total_sum + cache[504];
endrule
rule s506(sum_count == 506);
  total_sum <= total_sum + cache[505];
endrule
rule s507(sum_count == 507);
  total_sum <= total_sum + cache[506];
endrule
rule s508(sum_count == 508);
  total_sum <= total_sum + cache[507];
endrule
rule s509(sum_count == 509);
  total_sum <= total_sum + cache[508];
endrule
rule s510(sum_count == 510);
  total_sum <= total_sum + cache[509];
endrule
rule s511(sum_count == 511);
  total_sum <= total_sum + cache[510];
endrule
rule s512(sum_count == 512);
  total_sum <= total_sum + cache[511];
endrule
rule s513(sum_count == 513);
  total_sum <= total_sum + cache[512];
endrule
rule s514(sum_count == 514);
  total_sum <= total_sum + cache[513];
endrule
rule s515(sum_count == 515);
  total_sum <= total_sum + cache[514];
endrule
rule s516(sum_count == 516);
  total_sum <= total_sum + cache[515];
endrule
rule s517(sum_count == 517);
  total_sum <= total_sum + cache[516];
endrule
rule s518(sum_count == 518);
  total_sum <= total_sum + cache[517];
endrule
rule s519(sum_count == 519);
  total_sum <= total_sum + cache[518];
endrule
rule s520(sum_count == 520);
  total_sum <= total_sum + cache[519];
endrule
rule s521(sum_count == 521);
  total_sum <= total_sum + cache[520];
endrule
rule s522(sum_count == 522);
  total_sum <= total_sum + cache[521];
endrule
rule s523(sum_count == 523);
  total_sum <= total_sum + cache[522];
endrule
rule s524(sum_count == 524);
  total_sum <= total_sum + cache[523];
endrule
rule s525(sum_count == 525);
  total_sum <= total_sum + cache[524];
endrule
rule s526(sum_count == 526);
  total_sum <= total_sum + cache[525];
endrule
rule s527(sum_count == 527);
  total_sum <= total_sum + cache[526];
endrule
rule s528(sum_count == 528);
  total_sum <= total_sum + cache[527];
endrule
rule s529(sum_count == 529);
  total_sum <= total_sum + cache[528];
endrule
rule s530(sum_count == 530);
  total_sum <= total_sum + cache[529];
endrule
rule s531(sum_count == 531);
  total_sum <= total_sum + cache[530];
endrule
rule s532(sum_count == 532);
  total_sum <= total_sum + cache[531];
endrule
rule s533(sum_count == 533);
  total_sum <= total_sum + cache[532];
endrule
rule s534(sum_count == 534);
  total_sum <= total_sum + cache[533];
endrule
rule s535(sum_count == 535);
  total_sum <= total_sum + cache[534];
endrule
rule s536(sum_count == 536);
  total_sum <= total_sum + cache[535];
endrule
rule s537(sum_count == 537);
  total_sum <= total_sum + cache[536];
endrule
rule s538(sum_count == 538);
  total_sum <= total_sum + cache[537];
endrule
rule s539(sum_count == 539);
  total_sum <= total_sum + cache[538];
endrule
rule s540(sum_count == 540);
  total_sum <= total_sum + cache[539];
endrule
rule s541(sum_count == 541);
  total_sum <= total_sum + cache[540];
endrule
rule s542(sum_count == 542);
  total_sum <= total_sum + cache[541];
endrule
rule s543(sum_count == 543);
  total_sum <= total_sum + cache[542];
endrule
rule s544(sum_count == 544);
  total_sum <= total_sum + cache[543];
endrule
rule s545(sum_count == 545);
  total_sum <= total_sum + cache[544];
endrule
rule s546(sum_count == 546);
  total_sum <= total_sum + cache[545];
endrule
rule s547(sum_count == 547);
  total_sum <= total_sum + cache[546];
endrule
rule s548(sum_count == 548);
  total_sum <= total_sum + cache[547];
endrule
rule s549(sum_count == 549);
  total_sum <= total_sum + cache[548];
endrule
rule s550(sum_count == 550);
  total_sum <= total_sum + cache[549];
endrule
rule s551(sum_count == 551);
  total_sum <= total_sum + cache[550];
endrule
rule s552(sum_count == 552);
  total_sum <= total_sum + cache[551];
endrule
rule s553(sum_count == 553);
  total_sum <= total_sum + cache[552];
endrule
rule s554(sum_count == 554);
  total_sum <= total_sum + cache[553];
endrule
rule s555(sum_count == 555);
  total_sum <= total_sum + cache[554];
endrule
rule s556(sum_count == 556);
  total_sum <= total_sum + cache[555];
endrule
rule s557(sum_count == 557);
  total_sum <= total_sum + cache[556];
endrule
rule s558(sum_count == 558);
  total_sum <= total_sum + cache[557];
endrule
rule s559(sum_count == 559);
  total_sum <= total_sum + cache[558];
endrule
rule s560(sum_count == 560);
  total_sum <= total_sum + cache[559];
endrule
rule s561(sum_count == 561);
  total_sum <= total_sum + cache[560];
endrule
rule s562(sum_count == 562);
  total_sum <= total_sum + cache[561];
endrule
rule s563(sum_count == 563);
  total_sum <= total_sum + cache[562];
endrule
rule s564(sum_count == 564);
  total_sum <= total_sum + cache[563];
endrule
rule s565(sum_count == 565);
  total_sum <= total_sum + cache[564];
endrule
rule s566(sum_count == 566);
  total_sum <= total_sum + cache[565];
endrule
rule s567(sum_count == 567);
  total_sum <= total_sum + cache[566];
endrule
rule s568(sum_count == 568);
  total_sum <= total_sum + cache[567];
endrule
rule s569(sum_count == 569);
  total_sum <= total_sum + cache[568];
endrule
rule s570(sum_count == 570);
  total_sum <= total_sum + cache[569];
endrule
rule s571(sum_count == 571);
  total_sum <= total_sum + cache[570];
endrule
rule s572(sum_count == 572);
  total_sum <= total_sum + cache[571];
endrule
rule s573(sum_count == 573);
  total_sum <= total_sum + cache[572];
endrule
rule s574(sum_count == 574);
  total_sum <= total_sum + cache[573];
endrule
rule s575(sum_count == 575);
  total_sum <= total_sum + cache[574];
endrule
rule s576(sum_count == 576);
  total_sum <= total_sum + cache[575];
endrule
rule s577(sum_count == 577);
  total_sum <= total_sum + cache[576];
endrule
rule s578(sum_count == 578);
  total_sum <= total_sum + cache[577];
endrule
rule s579(sum_count == 579);
  total_sum <= total_sum + cache[578];
endrule
rule s580(sum_count == 580);
  total_sum <= total_sum + cache[579];
endrule
rule s581(sum_count == 581);
  total_sum <= total_sum + cache[580];
endrule
rule s582(sum_count == 582);
  total_sum <= total_sum + cache[581];
endrule
rule s583(sum_count == 583);
  total_sum <= total_sum + cache[582];
endrule
rule s584(sum_count == 584);
  total_sum <= total_sum + cache[583];
endrule
rule s585(sum_count == 585);
  total_sum <= total_sum + cache[584];
endrule
rule s586(sum_count == 586);
  total_sum <= total_sum + cache[585];
endrule
rule s587(sum_count == 587);
  total_sum <= total_sum + cache[586];
endrule
rule s588(sum_count == 588);
  total_sum <= total_sum + cache[587];
endrule
rule s589(sum_count == 589);
  total_sum <= total_sum + cache[588];
endrule
rule s590(sum_count == 590);
  total_sum <= total_sum + cache[589];
endrule
rule s591(sum_count == 591);
  total_sum <= total_sum + cache[590];
endrule
rule s592(sum_count == 592);
  total_sum <= total_sum + cache[591];
endrule
rule s593(sum_count == 593);
  total_sum <= total_sum + cache[592];
endrule
rule s594(sum_count == 594);
  total_sum <= total_sum + cache[593];
endrule
rule s595(sum_count == 595);
  total_sum <= total_sum + cache[594];
endrule
rule s596(sum_count == 596);
  total_sum <= total_sum + cache[595];
endrule
rule s597(sum_count == 597);
  total_sum <= total_sum + cache[596];
endrule
rule s598(sum_count == 598);
  total_sum <= total_sum + cache[597];
endrule
rule s599(sum_count == 599);
  total_sum <= total_sum + cache[598];
endrule
rule s600(sum_count == 600);
  total_sum <= total_sum + cache[599];
endrule
rule s601(sum_count == 601);
  total_sum <= total_sum + cache[600];
endrule
rule s602(sum_count == 602);
  total_sum <= total_sum + cache[601];
endrule
rule s603(sum_count == 603);
  total_sum <= total_sum + cache[602];
endrule
rule s604(sum_count == 604);
  total_sum <= total_sum + cache[603];
endrule
rule s605(sum_count == 605);
  total_sum <= total_sum + cache[604];
endrule
rule s606(sum_count == 606);
  total_sum <= total_sum + cache[605];
endrule
rule s607(sum_count == 607);
  total_sum <= total_sum + cache[606];
endrule
rule s608(sum_count == 608);
  total_sum <= total_sum + cache[607];
endrule
rule s609(sum_count == 609);
  total_sum <= total_sum + cache[608];
endrule
rule s610(sum_count == 610);
  total_sum <= total_sum + cache[609];
endrule
rule s611(sum_count == 611);
  total_sum <= total_sum + cache[610];
endrule
rule s612(sum_count == 612);
  total_sum <= total_sum + cache[611];
endrule
rule s613(sum_count == 613);
  total_sum <= total_sum + cache[612];
endrule
rule s614(sum_count == 614);
  total_sum <= total_sum + cache[613];
endrule
rule s615(sum_count == 615);
  total_sum <= total_sum + cache[614];
endrule
rule s616(sum_count == 616);
  total_sum <= total_sum + cache[615];
endrule
rule s617(sum_count == 617);
  total_sum <= total_sum + cache[616];
endrule
rule s618(sum_count == 618);
  total_sum <= total_sum + cache[617];
endrule
rule s619(sum_count == 619);
  total_sum <= total_sum + cache[618];
endrule
rule s620(sum_count == 620);
  total_sum <= total_sum + cache[619];
endrule
rule s621(sum_count == 621);
  total_sum <= total_sum + cache[620];
endrule
rule s622(sum_count == 622);
  total_sum <= total_sum + cache[621];
endrule
rule s623(sum_count == 623);
  total_sum <= total_sum + cache[622];
endrule
rule s624(sum_count == 624);
  total_sum <= total_sum + cache[623];
endrule
rule s625(sum_count == 625);
  total_sum <= total_sum + cache[624];
endrule
rule s626(sum_count == 626);
  total_sum <= total_sum + cache[625];
endrule
rule s627(sum_count == 627);
  total_sum <= total_sum + cache[626];
endrule
rule s628(sum_count == 628);
  total_sum <= total_sum + cache[627];
endrule
rule s629(sum_count == 629);
  total_sum <= total_sum + cache[628];
endrule
rule s630(sum_count == 630);
  total_sum <= total_sum + cache[629];
endrule
rule s631(sum_count == 631);
  total_sum <= total_sum + cache[630];
endrule
rule s632(sum_count == 632);
  total_sum <= total_sum + cache[631];
endrule
rule s633(sum_count == 633);
  total_sum <= total_sum + cache[632];
endrule
rule s634(sum_count == 634);
  total_sum <= total_sum + cache[633];
endrule
rule s635(sum_count == 635);
  total_sum <= total_sum + cache[634];
endrule
rule s636(sum_count == 636);
  total_sum <= total_sum + cache[635];
endrule
rule s637(sum_count == 637);
  total_sum <= total_sum + cache[636];
endrule
rule s638(sum_count == 638);
  total_sum <= total_sum + cache[637];
endrule
rule s639(sum_count == 639);
  total_sum <= total_sum + cache[638];
endrule
rule s640(sum_count == 640);
  total_sum <= total_sum + cache[639];
endrule
rule s641(sum_count == 641);
  total_sum <= total_sum + cache[640];
endrule
rule s642(sum_count == 642);
  total_sum <= total_sum + cache[641];
endrule
rule s643(sum_count == 643);
  total_sum <= total_sum + cache[642];
endrule
rule s644(sum_count == 644);
  total_sum <= total_sum + cache[643];
endrule
rule s645(sum_count == 645);
  total_sum <= total_sum + cache[644];
endrule
rule s646(sum_count == 646);
  total_sum <= total_sum + cache[645];
endrule
rule s647(sum_count == 647);
  total_sum <= total_sum + cache[646];
endrule
rule s648(sum_count == 648);
  total_sum <= total_sum + cache[647];
endrule
rule s649(sum_count == 649);
  total_sum <= total_sum + cache[648];
endrule
rule s650(sum_count == 650);
  total_sum <= total_sum + cache[649];
endrule
rule s651(sum_count == 651);
  total_sum <= total_sum + cache[650];
endrule
rule s652(sum_count == 652);
  total_sum <= total_sum + cache[651];
endrule
rule s653(sum_count == 653);
  total_sum <= total_sum + cache[652];
endrule
rule s654(sum_count == 654);
  total_sum <= total_sum + cache[653];
endrule
rule s655(sum_count == 655);
  total_sum <= total_sum + cache[654];
endrule
rule s656(sum_count == 656);
  total_sum <= total_sum + cache[655];
endrule
rule s657(sum_count == 657);
  total_sum <= total_sum + cache[656];
endrule
rule s658(sum_count == 658);
  total_sum <= total_sum + cache[657];
endrule
rule s659(sum_count == 659);
  total_sum <= total_sum + cache[658];
endrule
rule s660(sum_count == 660);
  total_sum <= total_sum + cache[659];
endrule
rule s661(sum_count == 661);
  total_sum <= total_sum + cache[660];
endrule
rule s662(sum_count == 662);
  total_sum <= total_sum + cache[661];
endrule
rule s663(sum_count == 663);
  total_sum <= total_sum + cache[662];
endrule
rule s664(sum_count == 664);
  total_sum <= total_sum + cache[663];
endrule
rule s665(sum_count == 665);
  total_sum <= total_sum + cache[664];
endrule
rule s666(sum_count == 666);
  total_sum <= total_sum + cache[665];
endrule
rule s667(sum_count == 667);
  total_sum <= total_sum + cache[666];
endrule
rule s668(sum_count == 668);
  total_sum <= total_sum + cache[667];
endrule
rule s669(sum_count == 669);
  total_sum <= total_sum + cache[668];
endrule
rule s670(sum_count == 670);
  total_sum <= total_sum + cache[669];
endrule
rule s671(sum_count == 671);
  total_sum <= total_sum + cache[670];
endrule
rule s672(sum_count == 672);
  total_sum <= total_sum + cache[671];
endrule
rule s673(sum_count == 673);
  total_sum <= total_sum + cache[672];
endrule
rule s674(sum_count == 674);
  total_sum <= total_sum + cache[673];
endrule
rule s675(sum_count == 675);
  total_sum <= total_sum + cache[674];
endrule
rule s676(sum_count == 676);
  total_sum <= total_sum + cache[675];
endrule
rule s677(sum_count == 677);
  total_sum <= total_sum + cache[676];
endrule
rule s678(sum_count == 678);
  total_sum <= total_sum + cache[677];
endrule
rule s679(sum_count == 679);
  total_sum <= total_sum + cache[678];
endrule
rule s680(sum_count == 680);
  total_sum <= total_sum + cache[679];
endrule
rule s681(sum_count == 681);
  total_sum <= total_sum + cache[680];
endrule
rule s682(sum_count == 682);
  total_sum <= total_sum + cache[681];
endrule
rule s683(sum_count == 683);
  total_sum <= total_sum + cache[682];
endrule
rule s684(sum_count == 684);
  total_sum <= total_sum + cache[683];
endrule
rule s685(sum_count == 685);
  total_sum <= total_sum + cache[684];
endrule
rule s686(sum_count == 686);
  total_sum <= total_sum + cache[685];
endrule
rule s687(sum_count == 687);
  total_sum <= total_sum + cache[686];
endrule
rule s688(sum_count == 688);
  total_sum <= total_sum + cache[687];
endrule
rule s689(sum_count == 689);
  total_sum <= total_sum + cache[688];
endrule
rule s690(sum_count == 690);
  total_sum <= total_sum + cache[689];
endrule
rule s691(sum_count == 691);
  total_sum <= total_sum + cache[690];
endrule
rule s692(sum_count == 692);
  total_sum <= total_sum + cache[691];
endrule
rule s693(sum_count == 693);
  total_sum <= total_sum + cache[692];
endrule
rule s694(sum_count == 694);
  total_sum <= total_sum + cache[693];
endrule
rule s695(sum_count == 695);
  total_sum <= total_sum + cache[694];
endrule
rule s696(sum_count == 696);
  total_sum <= total_sum + cache[695];
endrule
rule s697(sum_count == 697);
  total_sum <= total_sum + cache[696];
endrule
rule s698(sum_count == 698);
  total_sum <= total_sum + cache[697];
endrule
rule s699(sum_count == 699);
  total_sum <= total_sum + cache[698];
endrule
rule s700(sum_count == 700);
  total_sum <= total_sum + cache[699];
endrule
rule s701(sum_count == 701);
  total_sum <= total_sum + cache[700];
endrule
rule s702(sum_count == 702);
  total_sum <= total_sum + cache[701];
endrule
rule s703(sum_count == 703);
  total_sum <= total_sum + cache[702];
endrule
rule s704(sum_count == 704);
  total_sum <= total_sum + cache[703];
endrule
rule s705(sum_count == 705);
  total_sum <= total_sum + cache[704];
endrule
rule s706(sum_count == 706);
  total_sum <= total_sum + cache[705];
endrule
rule s707(sum_count == 707);
  total_sum <= total_sum + cache[706];
endrule
rule s708(sum_count == 708);
  total_sum <= total_sum + cache[707];
endrule
rule s709(sum_count == 709);
  total_sum <= total_sum + cache[708];
endrule
rule s710(sum_count == 710);
  total_sum <= total_sum + cache[709];
endrule
rule s711(sum_count == 711);
  total_sum <= total_sum + cache[710];
endrule
rule s712(sum_count == 712);
  total_sum <= total_sum + cache[711];
endrule
rule s713(sum_count == 713);
  total_sum <= total_sum + cache[712];
endrule
rule s714(sum_count == 714);
  total_sum <= total_sum + cache[713];
endrule
rule s715(sum_count == 715);
  total_sum <= total_sum + cache[714];
endrule
rule s716(sum_count == 716);
  total_sum <= total_sum + cache[715];
endrule
rule s717(sum_count == 717);
  total_sum <= total_sum + cache[716];
endrule
rule s718(sum_count == 718);
  total_sum <= total_sum + cache[717];
endrule
rule s719(sum_count == 719);
  total_sum <= total_sum + cache[718];
endrule
rule s720(sum_count == 720);
  total_sum <= total_sum + cache[719];
endrule
rule s721(sum_count == 721);
  total_sum <= total_sum + cache[720];
endrule
rule s722(sum_count == 722);
  total_sum <= total_sum + cache[721];
endrule
rule s723(sum_count == 723);
  total_sum <= total_sum + cache[722];
endrule
rule s724(sum_count == 724);
  total_sum <= total_sum + cache[723];
endrule
rule s725(sum_count == 725);
  total_sum <= total_sum + cache[724];
endrule
rule s726(sum_count == 726);
  total_sum <= total_sum + cache[725];
endrule
rule s727(sum_count == 727);
  total_sum <= total_sum + cache[726];
endrule
rule s728(sum_count == 728);
  total_sum <= total_sum + cache[727];
endrule
rule s729(sum_count == 729);
  total_sum <= total_sum + cache[728];
endrule
rule s730(sum_count == 730);
  total_sum <= total_sum + cache[729];
endrule
rule s731(sum_count == 731);
  total_sum <= total_sum + cache[730];
endrule
rule s732(sum_count == 732);
  total_sum <= total_sum + cache[731];
endrule
rule s733(sum_count == 733);
  total_sum <= total_sum + cache[732];
endrule
rule s734(sum_count == 734);
  total_sum <= total_sum + cache[733];
endrule
rule s735(sum_count == 735);
  total_sum <= total_sum + cache[734];
endrule
rule s736(sum_count == 736);
  total_sum <= total_sum + cache[735];
endrule
rule s737(sum_count == 737);
  total_sum <= total_sum + cache[736];
endrule
rule s738(sum_count == 738);
  total_sum <= total_sum + cache[737];
endrule
rule s739(sum_count == 739);
  total_sum <= total_sum + cache[738];
endrule
rule s740(sum_count == 740);
  total_sum <= total_sum + cache[739];
endrule
rule s741(sum_count == 741);
  total_sum <= total_sum + cache[740];
endrule
rule s742(sum_count == 742);
  total_sum <= total_sum + cache[741];
endrule
rule s743(sum_count == 743);
  total_sum <= total_sum + cache[742];
endrule
rule s744(sum_count == 744);
  total_sum <= total_sum + cache[743];
endrule
rule s745(sum_count == 745);
  total_sum <= total_sum + cache[744];
endrule
rule s746(sum_count == 746);
  total_sum <= total_sum + cache[745];
endrule
rule s747(sum_count == 747);
  total_sum <= total_sum + cache[746];
endrule
rule s748(sum_count == 748);
  total_sum <= total_sum + cache[747];
endrule
rule s749(sum_count == 749);
  total_sum <= total_sum + cache[748];
endrule
rule s750(sum_count == 750);
  total_sum <= total_sum + cache[749];
endrule
rule s751(sum_count == 751);
  total_sum <= total_sum + cache[750];
endrule
rule s752(sum_count == 752);
  total_sum <= total_sum + cache[751];
endrule
rule s753(sum_count == 753);
  total_sum <= total_sum + cache[752];
endrule
rule s754(sum_count == 754);
  total_sum <= total_sum + cache[753];
endrule
rule s755(sum_count == 755);
  total_sum <= total_sum + cache[754];
endrule
rule s756(sum_count == 756);
  total_sum <= total_sum + cache[755];
endrule
rule s757(sum_count == 757);
  total_sum <= total_sum + cache[756];
endrule
rule s758(sum_count == 758);
  total_sum <= total_sum + cache[757];
endrule
rule s759(sum_count == 759);
  total_sum <= total_sum + cache[758];
endrule
rule s760(sum_count == 760);
  total_sum <= total_sum + cache[759];
endrule
rule s761(sum_count == 761);
  total_sum <= total_sum + cache[760];
endrule
rule s762(sum_count == 762);
  total_sum <= total_sum + cache[761];
endrule
rule s763(sum_count == 763);
  total_sum <= total_sum + cache[762];
endrule
rule s764(sum_count == 764);
  total_sum <= total_sum + cache[763];
endrule
rule s765(sum_count == 765);
  total_sum <= total_sum + cache[764];
endrule
rule s766(sum_count == 766);
  total_sum <= total_sum + cache[765];
endrule
rule s767(sum_count == 767);
  total_sum <= total_sum + cache[766];
endrule
rule s768(sum_count == 768);
  total_sum <= total_sum + cache[767];
endrule
rule s769(sum_count == 769);
  total_sum <= total_sum + cache[768];
endrule
rule s770(sum_count == 770);
  total_sum <= total_sum + cache[769];
endrule
rule s771(sum_count == 771);
  total_sum <= total_sum + cache[770];
endrule
rule s772(sum_count == 772);
  total_sum <= total_sum + cache[771];
endrule
rule s773(sum_count == 773);
  total_sum <= total_sum + cache[772];
endrule
rule s774(sum_count == 774);
  total_sum <= total_sum + cache[773];
endrule
rule s775(sum_count == 775);
  total_sum <= total_sum + cache[774];
endrule
rule s776(sum_count == 776);
  total_sum <= total_sum + cache[775];
endrule
rule s777(sum_count == 777);
  total_sum <= total_sum + cache[776];
endrule
rule s778(sum_count == 778);
  total_sum <= total_sum + cache[777];
endrule
rule s779(sum_count == 779);
  total_sum <= total_sum + cache[778];
endrule
rule s780(sum_count == 780);
  total_sum <= total_sum + cache[779];
endrule
rule s781(sum_count == 781);
  total_sum <= total_sum + cache[780];
endrule
rule s782(sum_count == 782);
  total_sum <= total_sum + cache[781];
endrule
rule s783(sum_count == 783);
  total_sum <= total_sum + cache[782];
endrule
rule s784(sum_count == 784);
  total_sum <= total_sum + cache[783];
endrule
rule s785(sum_count == 785);
  total_sum <= total_sum + cache[784];
endrule
rule s786(sum_count == 786);
  total_sum <= total_sum + cache[785];
endrule
rule s787(sum_count == 787);
  total_sum <= total_sum + cache[786];
endrule
rule s788(sum_count == 788);
  total_sum <= total_sum + cache[787];
endrule
rule s789(sum_count == 789);
  total_sum <= total_sum + cache[788];
endrule
rule s790(sum_count == 790);
  total_sum <= total_sum + cache[789];
endrule
rule s791(sum_count == 791);
  total_sum <= total_sum + cache[790];
endrule
rule s792(sum_count == 792);
  total_sum <= total_sum + cache[791];
endrule
rule s793(sum_count == 793);
  total_sum <= total_sum + cache[792];
endrule
rule s794(sum_count == 794);
  total_sum <= total_sum + cache[793];
endrule
rule s795(sum_count == 795);
  total_sum <= total_sum + cache[794];
endrule
rule s796(sum_count == 796);
  total_sum <= total_sum + cache[795];
endrule
rule s797(sum_count == 797);
  total_sum <= total_sum + cache[796];
endrule
rule s798(sum_count == 798);
  total_sum <= total_sum + cache[797];
endrule
rule s799(sum_count == 799);
  total_sum <= total_sum + cache[798];
endrule
rule s800(sum_count == 800);
  total_sum <= total_sum + cache[799];
endrule
rule s801(sum_count == 801);
  total_sum <= total_sum + cache[800];
endrule
rule s802(sum_count == 802);
  total_sum <= total_sum + cache[801];
endrule
rule s803(sum_count == 803);
  total_sum <= total_sum + cache[802];
endrule
rule s804(sum_count == 804);
  total_sum <= total_sum + cache[803];
endrule
rule s805(sum_count == 805);
  total_sum <= total_sum + cache[804];
endrule
rule s806(sum_count == 806);
  total_sum <= total_sum + cache[805];
endrule
rule s807(sum_count == 807);
  total_sum <= total_sum + cache[806];
endrule
rule s808(sum_count == 808);
  total_sum <= total_sum + cache[807];
endrule
rule s809(sum_count == 809);
  total_sum <= total_sum + cache[808];
endrule
rule s810(sum_count == 810);
  total_sum <= total_sum + cache[809];
endrule
rule s811(sum_count == 811);
  total_sum <= total_sum + cache[810];
endrule
rule s812(sum_count == 812);
  total_sum <= total_sum + cache[811];
endrule
rule s813(sum_count == 813);
  total_sum <= total_sum + cache[812];
endrule
rule s814(sum_count == 814);
  total_sum <= total_sum + cache[813];
endrule
rule s815(sum_count == 815);
  total_sum <= total_sum + cache[814];
endrule
rule s816(sum_count == 816);
  total_sum <= total_sum + cache[815];
endrule
rule s817(sum_count == 817);
  total_sum <= total_sum + cache[816];
endrule
rule s818(sum_count == 818);
  total_sum <= total_sum + cache[817];
endrule
rule s819(sum_count == 819);
  total_sum <= total_sum + cache[818];
endrule
rule s820(sum_count == 820);
  total_sum <= total_sum + cache[819];
endrule
rule s821(sum_count == 821);
  total_sum <= total_sum + cache[820];
endrule
rule s822(sum_count == 822);
  total_sum <= total_sum + cache[821];
endrule
rule s823(sum_count == 823);
  total_sum <= total_sum + cache[822];
endrule
rule s824(sum_count == 824);
  total_sum <= total_sum + cache[823];
endrule
rule s825(sum_count == 825);
  total_sum <= total_sum + cache[824];
endrule
rule s826(sum_count == 826);
  total_sum <= total_sum + cache[825];
endrule
rule s827(sum_count == 827);
  total_sum <= total_sum + cache[826];
endrule
rule s828(sum_count == 828);
  total_sum <= total_sum + cache[827];
endrule
rule s829(sum_count == 829);
  total_sum <= total_sum + cache[828];
endrule
rule s830(sum_count == 830);
  total_sum <= total_sum + cache[829];
endrule
rule s831(sum_count == 831);
  total_sum <= total_sum + cache[830];
endrule
rule s832(sum_count == 832);
  total_sum <= total_sum + cache[831];
endrule
rule s833(sum_count == 833);
  total_sum <= total_sum + cache[832];
endrule
rule s834(sum_count == 834);
  total_sum <= total_sum + cache[833];
endrule
rule s835(sum_count == 835);
  total_sum <= total_sum + cache[834];
endrule
rule s836(sum_count == 836);
  total_sum <= total_sum + cache[835];
endrule
rule s837(sum_count == 837);
  total_sum <= total_sum + cache[836];
endrule
rule s838(sum_count == 838);
  total_sum <= total_sum + cache[837];
endrule
rule s839(sum_count == 839);
  total_sum <= total_sum + cache[838];
endrule
rule s840(sum_count == 840);
  total_sum <= total_sum + cache[839];
endrule
rule s841(sum_count == 841);
  total_sum <= total_sum + cache[840];
endrule
rule s842(sum_count == 842);
  total_sum <= total_sum + cache[841];
endrule
rule s843(sum_count == 843);
  total_sum <= total_sum + cache[842];
endrule
rule s844(sum_count == 844);
  total_sum <= total_sum + cache[843];
endrule
rule s845(sum_count == 845);
  total_sum <= total_sum + cache[844];
endrule
rule s846(sum_count == 846);
  total_sum <= total_sum + cache[845];
endrule
rule s847(sum_count == 847);
  total_sum <= total_sum + cache[846];
endrule
rule s848(sum_count == 848);
  total_sum <= total_sum + cache[847];
endrule
rule s849(sum_count == 849);
  total_sum <= total_sum + cache[848];
endrule
rule s850(sum_count == 850);
  total_sum <= total_sum + cache[849];
endrule
rule s851(sum_count == 851);
  total_sum <= total_sum + cache[850];
endrule
rule s852(sum_count == 852);
  total_sum <= total_sum + cache[851];
endrule
rule s853(sum_count == 853);
  total_sum <= total_sum + cache[852];
endrule
rule s854(sum_count == 854);
  total_sum <= total_sum + cache[853];
endrule
rule s855(sum_count == 855);
  total_sum <= total_sum + cache[854];
endrule
rule s856(sum_count == 856);
  total_sum <= total_sum + cache[855];
endrule
rule s857(sum_count == 857);
  total_sum <= total_sum + cache[856];
endrule
rule s858(sum_count == 858);
  total_sum <= total_sum + cache[857];
endrule
rule s859(sum_count == 859);
  total_sum <= total_sum + cache[858];
endrule
rule s860(sum_count == 860);
  total_sum <= total_sum + cache[859];
endrule
rule s861(sum_count == 861);
  total_sum <= total_sum + cache[860];
endrule
rule s862(sum_count == 862);
  total_sum <= total_sum + cache[861];
endrule
rule s863(sum_count == 863);
  total_sum <= total_sum + cache[862];
endrule
rule s864(sum_count == 864);
  total_sum <= total_sum + cache[863];
endrule
rule s865(sum_count == 865);
  total_sum <= total_sum + cache[864];
endrule
rule s866(sum_count == 866);
  total_sum <= total_sum + cache[865];
endrule
rule s867(sum_count == 867);
  total_sum <= total_sum + cache[866];
endrule
rule s868(sum_count == 868);
  total_sum <= total_sum + cache[867];
endrule
rule s869(sum_count == 869);
  total_sum <= total_sum + cache[868];
endrule
rule s870(sum_count == 870);
  total_sum <= total_sum + cache[869];
endrule
rule s871(sum_count == 871);
  total_sum <= total_sum + cache[870];
endrule
rule s872(sum_count == 872);
  total_sum <= total_sum + cache[871];
endrule
rule s873(sum_count == 873);
  total_sum <= total_sum + cache[872];
endrule
rule s874(sum_count == 874);
  total_sum <= total_sum + cache[873];
endrule
rule s875(sum_count == 875);
  total_sum <= total_sum + cache[874];
endrule
rule s876(sum_count == 876);
  total_sum <= total_sum + cache[875];
endrule
rule s877(sum_count == 877);
  total_sum <= total_sum + cache[876];
endrule
rule s878(sum_count == 878);
  total_sum <= total_sum + cache[877];
endrule
rule s879(sum_count == 879);
  total_sum <= total_sum + cache[878];
endrule
rule s880(sum_count == 880);
  total_sum <= total_sum + cache[879];
endrule
rule s881(sum_count == 881);
  total_sum <= total_sum + cache[880];
endrule
rule s882(sum_count == 882);
  total_sum <= total_sum + cache[881];
endrule
rule s883(sum_count == 883);
  total_sum <= total_sum + cache[882];
endrule
rule s884(sum_count == 884);
  total_sum <= total_sum + cache[883];
endrule
rule s885(sum_count == 885);
  total_sum <= total_sum + cache[884];
endrule
rule s886(sum_count == 886);
  total_sum <= total_sum + cache[885];
endrule
rule s887(sum_count == 887);
  total_sum <= total_sum + cache[886];
endrule
rule s888(sum_count == 888);
  total_sum <= total_sum + cache[887];
endrule
rule s889(sum_count == 889);
  total_sum <= total_sum + cache[888];
endrule
rule s890(sum_count == 890);
  total_sum <= total_sum + cache[889];
endrule
rule s891(sum_count == 891);
  total_sum <= total_sum + cache[890];
endrule
rule s892(sum_count == 892);
  total_sum <= total_sum + cache[891];
endrule
rule s893(sum_count == 893);
  total_sum <= total_sum + cache[892];
endrule
rule s894(sum_count == 894);
  total_sum <= total_sum + cache[893];
endrule
rule s895(sum_count == 895);
  total_sum <= total_sum + cache[894];
endrule
rule s896(sum_count == 896);
  total_sum <= total_sum + cache[895];
endrule
rule s897(sum_count == 897);
  total_sum <= total_sum + cache[896];
endrule
rule s898(sum_count == 898);
  total_sum <= total_sum + cache[897];
endrule
rule s899(sum_count == 899);
  total_sum <= total_sum + cache[898];
endrule
rule s900(sum_count == 900);
  total_sum <= total_sum + cache[899];
endrule
rule s901(sum_count == 901);
  total_sum <= total_sum + cache[900];
endrule
rule s902(sum_count == 902);
  total_sum <= total_sum + cache[901];
endrule
rule s903(sum_count == 903);
  total_sum <= total_sum + cache[902];
endrule
rule s904(sum_count == 904);
  total_sum <= total_sum + cache[903];
endrule
rule s905(sum_count == 905);
  total_sum <= total_sum + cache[904];
endrule
rule s906(sum_count == 906);
  total_sum <= total_sum + cache[905];
endrule
rule s907(sum_count == 907);
  total_sum <= total_sum + cache[906];
endrule
rule s908(sum_count == 908);
  total_sum <= total_sum + cache[907];
endrule
rule s909(sum_count == 909);
  total_sum <= total_sum + cache[908];
endrule
rule s910(sum_count == 910);
  total_sum <= total_sum + cache[909];
endrule
rule s911(sum_count == 911);
  total_sum <= total_sum + cache[910];
endrule
rule s912(sum_count == 912);
  total_sum <= total_sum + cache[911];
endrule
rule s913(sum_count == 913);
  total_sum <= total_sum + cache[912];
endrule
rule s914(sum_count == 914);
  total_sum <= total_sum + cache[913];
endrule
rule s915(sum_count == 915);
  total_sum <= total_sum + cache[914];
endrule
rule s916(sum_count == 916);
  total_sum <= total_sum + cache[915];
endrule
rule s917(sum_count == 917);
  total_sum <= total_sum + cache[916];
endrule
rule s918(sum_count == 918);
  total_sum <= total_sum + cache[917];
endrule
rule s919(sum_count == 919);
  total_sum <= total_sum + cache[918];
endrule
rule s920(sum_count == 920);
  total_sum <= total_sum + cache[919];
endrule
rule s921(sum_count == 921);
  total_sum <= total_sum + cache[920];
endrule
rule s922(sum_count == 922);
  total_sum <= total_sum + cache[921];
endrule
rule s923(sum_count == 923);
  total_sum <= total_sum + cache[922];
endrule
rule s924(sum_count == 924);
  total_sum <= total_sum + cache[923];
endrule
rule s925(sum_count == 925);
  total_sum <= total_sum + cache[924];
endrule
rule s926(sum_count == 926);
  total_sum <= total_sum + cache[925];
endrule
rule s927(sum_count == 927);
  total_sum <= total_sum + cache[926];
endrule
rule s928(sum_count == 928);
  total_sum <= total_sum + cache[927];
endrule
rule s929(sum_count == 929);
  total_sum <= total_sum + cache[928];
endrule
rule s930(sum_count == 930);
  total_sum <= total_sum + cache[929];
endrule
rule s931(sum_count == 931);
  total_sum <= total_sum + cache[930];
endrule
rule s932(sum_count == 932);
  total_sum <= total_sum + cache[931];
endrule
rule s933(sum_count == 933);
  total_sum <= total_sum + cache[932];
endrule
rule s934(sum_count == 934);
  total_sum <= total_sum + cache[933];
endrule
rule s935(sum_count == 935);
  total_sum <= total_sum + cache[934];
endrule
rule s936(sum_count == 936);
  total_sum <= total_sum + cache[935];
endrule
rule s937(sum_count == 937);
  total_sum <= total_sum + cache[936];
endrule
rule s938(sum_count == 938);
  total_sum <= total_sum + cache[937];
endrule
rule s939(sum_count == 939);
  total_sum <= total_sum + cache[938];
endrule
rule s940(sum_count == 940);
  total_sum <= total_sum + cache[939];
endrule
rule s941(sum_count == 941);
  total_sum <= total_sum + cache[940];
endrule
rule s942(sum_count == 942);
  total_sum <= total_sum + cache[941];
endrule
rule s943(sum_count == 943);
  total_sum <= total_sum + cache[942];
endrule
rule s944(sum_count == 944);
  total_sum <= total_sum + cache[943];
endrule
rule s945(sum_count == 945);
  total_sum <= total_sum + cache[944];
endrule
rule s946(sum_count == 946);
  total_sum <= total_sum + cache[945];
endrule
rule s947(sum_count == 947);
  total_sum <= total_sum + cache[946];
endrule
rule s948(sum_count == 948);
  total_sum <= total_sum + cache[947];
endrule
rule s949(sum_count == 949);
  total_sum <= total_sum + cache[948];
endrule
rule s950(sum_count == 950);
  total_sum <= total_sum + cache[949];
endrule
rule s951(sum_count == 951);
  total_sum <= total_sum + cache[950];
endrule
rule s952(sum_count == 952);
  total_sum <= total_sum + cache[951];
endrule
rule s953(sum_count == 953);
  total_sum <= total_sum + cache[952];
endrule
rule s954(sum_count == 954);
  total_sum <= total_sum + cache[953];
endrule
rule s955(sum_count == 955);
  total_sum <= total_sum + cache[954];
endrule
rule s956(sum_count == 956);
  total_sum <= total_sum + cache[955];
endrule
rule s957(sum_count == 957);
  total_sum <= total_sum + cache[956];
endrule
rule s958(sum_count == 958);
  total_sum <= total_sum + cache[957];
endrule
rule s959(sum_count == 959);
  total_sum <= total_sum + cache[958];
endrule
rule s960(sum_count == 960);
  total_sum <= total_sum + cache[959];
endrule
rule s961(sum_count == 961);
  total_sum <= total_sum + cache[960];
endrule
rule s962(sum_count == 962);
  total_sum <= total_sum + cache[961];
endrule
rule s963(sum_count == 963);
  total_sum <= total_sum + cache[962];
endrule
rule s964(sum_count == 964);
  total_sum <= total_sum + cache[963];
endrule
rule s965(sum_count == 965);
  total_sum <= total_sum + cache[964];
endrule
rule s966(sum_count == 966);
  total_sum <= total_sum + cache[965];
endrule
rule s967(sum_count == 967);
  total_sum <= total_sum + cache[966];
endrule
rule s968(sum_count == 968);
  total_sum <= total_sum + cache[967];
endrule
rule s969(sum_count == 969);
  total_sum <= total_sum + cache[968];
endrule
rule s970(sum_count == 970);
  total_sum <= total_sum + cache[969];
endrule
rule s971(sum_count == 971);
  total_sum <= total_sum + cache[970];
endrule
rule s972(sum_count == 972);
  total_sum <= total_sum + cache[971];
endrule
rule s973(sum_count == 973);
  total_sum <= total_sum + cache[972];
endrule
rule s974(sum_count == 974);
  total_sum <= total_sum + cache[973];
endrule
rule s975(sum_count == 975);
  total_sum <= total_sum + cache[974];
endrule
rule s976(sum_count == 976);
  total_sum <= total_sum + cache[975];
endrule
rule s977(sum_count == 977);
  total_sum <= total_sum + cache[976];
endrule
rule s978(sum_count == 978);
  total_sum <= total_sum + cache[977];
endrule
rule s979(sum_count == 979);
  total_sum <= total_sum + cache[978];
endrule
rule s980(sum_count == 980);
  total_sum <= total_sum + cache[979];
endrule
rule s981(sum_count == 981);
  total_sum <= total_sum + cache[980];
endrule
rule s982(sum_count == 982);
  total_sum <= total_sum + cache[981];
endrule
rule s983(sum_count == 983);
  total_sum <= total_sum + cache[982];
endrule
rule s984(sum_count == 984);
  total_sum <= total_sum + cache[983];
endrule
rule s985(sum_count == 985);
  total_sum <= total_sum + cache[984];
endrule
rule s986(sum_count == 986);
  total_sum <= total_sum + cache[985];
endrule
rule s987(sum_count == 987);
  total_sum <= total_sum + cache[986];
endrule
rule s988(sum_count == 988);
  total_sum <= total_sum + cache[987];
endrule
rule s989(sum_count == 989);
  total_sum <= total_sum + cache[988];
endrule
rule s990(sum_count == 990);
  total_sum <= total_sum + cache[989];
endrule
rule s991(sum_count == 991);
  total_sum <= total_sum + cache[990];
endrule
rule s992(sum_count == 992);
  total_sum <= total_sum + cache[991];
endrule
rule s993(sum_count == 993);
  total_sum <= total_sum + cache[992];
endrule
rule s994(sum_count == 994);
  total_sum <= total_sum + cache[993];
endrule
rule s995(sum_count == 995);
  total_sum <= total_sum + cache[994];
endrule
rule s996(sum_count == 996);
  total_sum <= total_sum + cache[995];
endrule
rule s997(sum_count == 997);
  total_sum <= total_sum + cache[996];
endrule
rule s998(sum_count == 998);
  total_sum <= total_sum + cache[997];
endrule
rule s999(sum_count == 999);
  total_sum <= total_sum + cache[998];
endrule
rule s1000(sum_count == 1000);
  total_sum <= total_sum + cache[999];
endrule
rule s1001(sum_count == 1001);
  total_sum <= total_sum + cache[1000];
endrule
rule s1002(sum_count == 1002);
  total_sum <= total_sum + cache[1001];
endrule
rule s1003(sum_count == 1003);
  total_sum <= total_sum + cache[1002];
endrule
rule s1004(sum_count == 1004);
  total_sum <= total_sum + cache[1003];
endrule
rule s1005(sum_count == 1005);
  total_sum <= total_sum + cache[1004];
endrule
rule s1006(sum_count == 1006);
  total_sum <= total_sum + cache[1005];
endrule
rule s1007(sum_count == 1007);
  total_sum <= total_sum + cache[1006];
endrule
rule s1008(sum_count == 1008);
  total_sum <= total_sum + cache[1007];
endrule
rule s1009(sum_count == 1009);
  total_sum <= total_sum + cache[1008];
endrule
rule s1010(sum_count == 1010);
  total_sum <= total_sum + cache[1009];
endrule
rule s1011(sum_count == 1011);
  total_sum <= total_sum + cache[1010];
endrule
rule s1012(sum_count == 1012);
  total_sum <= total_sum + cache[1011];
endrule
rule s1013(sum_count == 1013);
  total_sum <= total_sum + cache[1012];
endrule
rule s1014(sum_count == 1014);
  total_sum <= total_sum + cache[1013];
endrule
rule s1015(sum_count == 1015);
  total_sum <= total_sum + cache[1014];
endrule
rule s1016(sum_count == 1016);
  total_sum <= total_sum + cache[1015];
endrule
rule s1017(sum_count == 1017);
  total_sum <= total_sum + cache[1016];
endrule
rule s1018(sum_count == 1018);
  total_sum <= total_sum + cache[1017];
endrule
rule s1019(sum_count == 1019);
  total_sum <= total_sum + cache[1018];
endrule
rule s1020(sum_count == 1020);
  total_sum <= total_sum + cache[1019];
endrule
rule s1021(sum_count == 1021);
  total_sum <= total_sum + cache[1020];
endrule
rule s1022(sum_count == 1022);
  total_sum <= total_sum + cache[1021];
endrule
rule s1023(sum_count == 1023);
  total_sum <= total_sum + cache[1022];
endrule
rule s1024(sum_count == 1024);
  total_sum <= total_sum + cache[1023];
endrule
rule s1025(sum_count == 1025);
  total_sum <= total_sum + cache[1024];
endrule
rule s1026(sum_count == 1026);
  total_sum <= total_sum + cache[1025];
endrule
rule s1027(sum_count == 1027);
  total_sum <= total_sum + cache[1026];
endrule
rule s1028(sum_count == 1028);
  total_sum <= total_sum + cache[1027];
endrule
rule s1029(sum_count == 1029);
  total_sum <= total_sum + cache[1028];
endrule
rule s1030(sum_count == 1030);
  total_sum <= total_sum + cache[1029];
endrule
rule s1031(sum_count == 1031);
  total_sum <= total_sum + cache[1030];
endrule
rule s1032(sum_count == 1032);
  total_sum <= total_sum + cache[1031];
endrule
rule s1033(sum_count == 1033);
  total_sum <= total_sum + cache[1032];
endrule
rule s1034(sum_count == 1034);
  total_sum <= total_sum + cache[1033];
endrule
rule s1035(sum_count == 1035);
  total_sum <= total_sum + cache[1034];
endrule
rule s1036(sum_count == 1036);
  total_sum <= total_sum + cache[1035];
endrule
rule s1037(sum_count == 1037);
  total_sum <= total_sum + cache[1036];
endrule
rule s1038(sum_count == 1038);
  total_sum <= total_sum + cache[1037];
endrule
rule s1039(sum_count == 1039);
  total_sum <= total_sum + cache[1038];
endrule
rule s1040(sum_count == 1040);
  total_sum <= total_sum + cache[1039];
endrule
rule s1041(sum_count == 1041);
  total_sum <= total_sum + cache[1040];
endrule
rule s1042(sum_count == 1042);
  total_sum <= total_sum + cache[1041];
endrule
rule s1043(sum_count == 1043);
  total_sum <= total_sum + cache[1042];
endrule
rule s1044(sum_count == 1044);
  total_sum <= total_sum + cache[1043];
endrule
rule s1045(sum_count == 1045);
  total_sum <= total_sum + cache[1044];
endrule
rule s1046(sum_count == 1046);
  total_sum <= total_sum + cache[1045];
endrule
rule s1047(sum_count == 1047);
  total_sum <= total_sum + cache[1046];
endrule
rule s1048(sum_count == 1048);
  total_sum <= total_sum + cache[1047];
endrule
rule s1049(sum_count == 1049);
  total_sum <= total_sum + cache[1048];
endrule
rule s1050(sum_count == 1050);
  total_sum <= total_sum + cache[1049];
endrule
rule s1051(sum_count == 1051);
  total_sum <= total_sum + cache[1050];
endrule
rule s1052(sum_count == 1052);
  total_sum <= total_sum + cache[1051];
endrule
rule s1053(sum_count == 1053);
  total_sum <= total_sum + cache[1052];
endrule
rule s1054(sum_count == 1054);
  total_sum <= total_sum + cache[1053];
endrule
rule s1055(sum_count == 1055);
  total_sum <= total_sum + cache[1054];
endrule
rule s1056(sum_count == 1056);
  total_sum <= total_sum + cache[1055];
endrule
rule s1057(sum_count == 1057);
  total_sum <= total_sum + cache[1056];
endrule
rule s1058(sum_count == 1058);
  total_sum <= total_sum + cache[1057];
endrule
rule s1059(sum_count == 1059);
  total_sum <= total_sum + cache[1058];
endrule
rule s1060(sum_count == 1060);
  total_sum <= total_sum + cache[1059];
endrule
rule s1061(sum_count == 1061);
  total_sum <= total_sum + cache[1060];
endrule
rule s1062(sum_count == 1062);
  total_sum <= total_sum + cache[1061];
endrule
rule s1063(sum_count == 1063);
  total_sum <= total_sum + cache[1062];
endrule
rule s1064(sum_count == 1064);
  total_sum <= total_sum + cache[1063];
endrule
rule s1065(sum_count == 1065);
  total_sum <= total_sum + cache[1064];
endrule
rule s1066(sum_count == 1066);
  total_sum <= total_sum + cache[1065];
endrule
rule s1067(sum_count == 1067);
  total_sum <= total_sum + cache[1066];
endrule
rule s1068(sum_count == 1068);
  total_sum <= total_sum + cache[1067];
endrule
rule s1069(sum_count == 1069);
  total_sum <= total_sum + cache[1068];
endrule
rule s1070(sum_count == 1070);
  total_sum <= total_sum + cache[1069];
endrule
rule s1071(sum_count == 1071);
  total_sum <= total_sum + cache[1070];
endrule
rule s1072(sum_count == 1072);
  total_sum <= total_sum + cache[1071];
endrule
rule s1073(sum_count == 1073);
  total_sum <= total_sum + cache[1072];
endrule
rule s1074(sum_count == 1074);
  total_sum <= total_sum + cache[1073];
endrule
rule s1075(sum_count == 1075);
  total_sum <= total_sum + cache[1074];
endrule
rule s1076(sum_count == 1076);
  total_sum <= total_sum + cache[1075];
endrule
rule s1077(sum_count == 1077);
  total_sum <= total_sum + cache[1076];
endrule
rule s1078(sum_count == 1078);
  total_sum <= total_sum + cache[1077];
endrule
rule s1079(sum_count == 1079);
  total_sum <= total_sum + cache[1078];
endrule
rule s1080(sum_count == 1080);
  total_sum <= total_sum + cache[1079];
endrule
rule s1081(sum_count == 1081);
  total_sum <= total_sum + cache[1080];
endrule
rule s1082(sum_count == 1082);
  total_sum <= total_sum + cache[1081];
endrule
rule s1083(sum_count == 1083);
  total_sum <= total_sum + cache[1082];
endrule
rule s1084(sum_count == 1084);
  total_sum <= total_sum + cache[1083];
endrule
rule s1085(sum_count == 1085);
  total_sum <= total_sum + cache[1084];
endrule
rule s1086(sum_count == 1086);
  total_sum <= total_sum + cache[1085];
endrule
rule s1087(sum_count == 1087);
  total_sum <= total_sum + cache[1086];
endrule
rule s1088(sum_count == 1088);
  total_sum <= total_sum + cache[1087];
endrule
rule s1089(sum_count == 1089);
  total_sum <= total_sum + cache[1088];
endrule
rule s1090(sum_count == 1090);
  total_sum <= total_sum + cache[1089];
endrule
rule s1091(sum_count == 1091);
  total_sum <= total_sum + cache[1090];
endrule
rule s1092(sum_count == 1092);
  total_sum <= total_sum + cache[1091];
endrule
rule s1093(sum_count == 1093);
  total_sum <= total_sum + cache[1092];
endrule
rule s1094(sum_count == 1094);
  total_sum <= total_sum + cache[1093];
endrule
rule s1095(sum_count == 1095);
  total_sum <= total_sum + cache[1094];
endrule
rule s1096(sum_count == 1096);
  total_sum <= total_sum + cache[1095];
endrule
rule s1097(sum_count == 1097);
  total_sum <= total_sum + cache[1096];
endrule
rule s1098(sum_count == 1098);
  total_sum <= total_sum + cache[1097];
endrule
rule s1099(sum_count == 1099);
  total_sum <= total_sum + cache[1098];
endrule
rule s1100(sum_count == 1100);
  total_sum <= total_sum + cache[1099];
endrule
rule s1101(sum_count == 1101);
  total_sum <= total_sum + cache[1100];
endrule
rule s1102(sum_count == 1102);
  total_sum <= total_sum + cache[1101];
endrule
rule s1103(sum_count == 1103);
  total_sum <= total_sum + cache[1102];
endrule
rule s1104(sum_count == 1104);
  total_sum <= total_sum + cache[1103];
endrule
rule s1105(sum_count == 1105);
  total_sum <= total_sum + cache[1104];
endrule
rule s1106(sum_count == 1106);
  total_sum <= total_sum + cache[1105];
endrule
rule s1107(sum_count == 1107);
  total_sum <= total_sum + cache[1106];
endrule
rule s1108(sum_count == 1108);
  total_sum <= total_sum + cache[1107];
endrule
rule s1109(sum_count == 1109);
  total_sum <= total_sum + cache[1108];
endrule
rule s1110(sum_count == 1110);
  total_sum <= total_sum + cache[1109];
endrule
rule s1111(sum_count == 1111);
  total_sum <= total_sum + cache[1110];
endrule
rule s1112(sum_count == 1112);
  total_sum <= total_sum + cache[1111];
endrule
rule s1113(sum_count == 1113);
  total_sum <= total_sum + cache[1112];
endrule
rule s1114(sum_count == 1114);
  total_sum <= total_sum + cache[1113];
endrule
rule s1115(sum_count == 1115);
  total_sum <= total_sum + cache[1114];
endrule
rule s1116(sum_count == 1116);
  total_sum <= total_sum + cache[1115];
endrule
rule s1117(sum_count == 1117);
  total_sum <= total_sum + cache[1116];
endrule
rule s1118(sum_count == 1118);
  total_sum <= total_sum + cache[1117];
endrule
rule s1119(sum_count == 1119);
  total_sum <= total_sum + cache[1118];
endrule
rule s1120(sum_count == 1120);
  total_sum <= total_sum + cache[1119];
endrule
rule s1121(sum_count == 1121);
  total_sum <= total_sum + cache[1120];
endrule
rule s1122(sum_count == 1122);
  total_sum <= total_sum + cache[1121];
endrule
rule s1123(sum_count == 1123);
  total_sum <= total_sum + cache[1122];
endrule
rule s1124(sum_count == 1124);
  total_sum <= total_sum + cache[1123];
endrule
rule s1125(sum_count == 1125);
  total_sum <= total_sum + cache[1124];
endrule
rule s1126(sum_count == 1126);
  total_sum <= total_sum + cache[1125];
endrule
rule s1127(sum_count == 1127);
  total_sum <= total_sum + cache[1126];
endrule
rule s1128(sum_count == 1128);
  total_sum <= total_sum + cache[1127];
endrule
rule s1129(sum_count == 1129);
  total_sum <= total_sum + cache[1128];
endrule
rule s1130(sum_count == 1130);
  total_sum <= total_sum + cache[1129];
endrule
rule s1131(sum_count == 1131);
  total_sum <= total_sum + cache[1130];
endrule
rule s1132(sum_count == 1132);
  total_sum <= total_sum + cache[1131];
endrule
rule s1133(sum_count == 1133);
  total_sum <= total_sum + cache[1132];
endrule
rule s1134(sum_count == 1134);
  total_sum <= total_sum + cache[1133];
endrule
rule s1135(sum_count == 1135);
  total_sum <= total_sum + cache[1134];
endrule
rule s1136(sum_count == 1136);
  total_sum <= total_sum + cache[1135];
endrule
rule s1137(sum_count == 1137);
  total_sum <= total_sum + cache[1136];
endrule
rule s1138(sum_count == 1138);
  total_sum <= total_sum + cache[1137];
endrule
rule s1139(sum_count == 1139);
  total_sum <= total_sum + cache[1138];
endrule
rule s1140(sum_count == 1140);
  total_sum <= total_sum + cache[1139];
endrule
rule s1141(sum_count == 1141);
  total_sum <= total_sum + cache[1140];
endrule
rule s1142(sum_count == 1142);
  total_sum <= total_sum + cache[1141];
endrule
rule s1143(sum_count == 1143);
  total_sum <= total_sum + cache[1142];
endrule
rule s1144(sum_count == 1144);
  total_sum <= total_sum + cache[1143];
endrule
rule s1145(sum_count == 1145);
  total_sum <= total_sum + cache[1144];
endrule
rule s1146(sum_count == 1146);
  total_sum <= total_sum + cache[1145];
endrule
rule s1147(sum_count == 1147);
  total_sum <= total_sum + cache[1146];
endrule
rule s1148(sum_count == 1148);
  total_sum <= total_sum + cache[1147];
endrule
rule s1149(sum_count == 1149);
  total_sum <= total_sum + cache[1148];
endrule
rule s1150(sum_count == 1150);
  total_sum <= total_sum + cache[1149];
endrule
rule s1151(sum_count == 1151);
  total_sum <= total_sum + cache[1150];
endrule
rule s1152(sum_count == 1152);
  total_sum <= total_sum + cache[1151];
endrule
rule s1153(sum_count == 1153);
  total_sum <= total_sum + cache[1152];
endrule
rule s1154(sum_count == 1154);
  total_sum <= total_sum + cache[1153];
endrule
rule s1155(sum_count == 1155);
  total_sum <= total_sum + cache[1154];
endrule
rule s1156(sum_count == 1156);
  total_sum <= total_sum + cache[1155];
endrule
rule s1157(sum_count == 1157);
  total_sum <= total_sum + cache[1156];
endrule
rule s1158(sum_count == 1158);
  total_sum <= total_sum + cache[1157];
endrule
rule s1159(sum_count == 1159);
  total_sum <= total_sum + cache[1158];
endrule
rule s1160(sum_count == 1160);
  total_sum <= total_sum + cache[1159];
endrule
rule s1161(sum_count == 1161);
  total_sum <= total_sum + cache[1160];
endrule
rule s1162(sum_count == 1162);
  total_sum <= total_sum + cache[1161];
endrule
rule s1163(sum_count == 1163);
  total_sum <= total_sum + cache[1162];
endrule
rule s1164(sum_count == 1164);
  total_sum <= total_sum + cache[1163];
endrule
rule s1165(sum_count == 1165);
  total_sum <= total_sum + cache[1164];
endrule
rule s1166(sum_count == 1166);
  total_sum <= total_sum + cache[1165];
endrule
rule s1167(sum_count == 1167);
  total_sum <= total_sum + cache[1166];
endrule
rule s1168(sum_count == 1168);
  total_sum <= total_sum + cache[1167];
endrule
rule s1169(sum_count == 1169);
  total_sum <= total_sum + cache[1168];
endrule
rule s1170(sum_count == 1170);
  total_sum <= total_sum + cache[1169];
endrule
rule s1171(sum_count == 1171);
  total_sum <= total_sum + cache[1170];
endrule
rule s1172(sum_count == 1172);
  total_sum <= total_sum + cache[1171];
endrule
rule s1173(sum_count == 1173);
  total_sum <= total_sum + cache[1172];
endrule
rule s1174(sum_count == 1174);
  total_sum <= total_sum + cache[1173];
endrule
rule s1175(sum_count == 1175);
  total_sum <= total_sum + cache[1174];
endrule
rule s1176(sum_count == 1176);
  total_sum <= total_sum + cache[1175];
endrule
rule s1177(sum_count == 1177);
  total_sum <= total_sum + cache[1176];
endrule
rule s1178(sum_count == 1178);
  total_sum <= total_sum + cache[1177];
endrule
rule s1179(sum_count == 1179);
  total_sum <= total_sum + cache[1178];
endrule
rule s1180(sum_count == 1180);
  total_sum <= total_sum + cache[1179];
endrule
rule s1181(sum_count == 1181);
  total_sum <= total_sum + cache[1180];
endrule
rule s1182(sum_count == 1182);
  total_sum <= total_sum + cache[1181];
endrule
rule s1183(sum_count == 1183);
  total_sum <= total_sum + cache[1182];
endrule
rule s1184(sum_count == 1184);
  total_sum <= total_sum + cache[1183];
endrule
rule s1185(sum_count == 1185);
  total_sum <= total_sum + cache[1184];
endrule
rule s1186(sum_count == 1186);
  total_sum <= total_sum + cache[1185];
endrule
rule s1187(sum_count == 1187);
  total_sum <= total_sum + cache[1186];
endrule
rule s1188(sum_count == 1188);
  total_sum <= total_sum + cache[1187];
endrule
rule s1189(sum_count == 1189);
  total_sum <= total_sum + cache[1188];
endrule
rule s1190(sum_count == 1190);
  total_sum <= total_sum + cache[1189];
endrule
rule s1191(sum_count == 1191);
  total_sum <= total_sum + cache[1190];
endrule
rule s1192(sum_count == 1192);
  total_sum <= total_sum + cache[1191];
endrule
rule s1193(sum_count == 1193);
  total_sum <= total_sum + cache[1192];
endrule
rule s1194(sum_count == 1194);
  total_sum <= total_sum + cache[1193];
endrule
rule s1195(sum_count == 1195);
  total_sum <= total_sum + cache[1194];
endrule
rule s1196(sum_count == 1196);
  total_sum <= total_sum + cache[1195];
endrule
rule s1197(sum_count == 1197);
  total_sum <= total_sum + cache[1196];
endrule
rule s1198(sum_count == 1198);
  total_sum <= total_sum + cache[1197];
endrule
rule s1199(sum_count == 1199);
  total_sum <= total_sum + cache[1198];
endrule
rule s1200(sum_count == 1200);
  total_sum <= total_sum + cache[1199];
endrule
rule s1201(sum_count == 1201);
  total_sum <= total_sum + cache[1200];
endrule
rule s1202(sum_count == 1202);
  total_sum <= total_sum + cache[1201];
endrule
rule s1203(sum_count == 1203);
  total_sum <= total_sum + cache[1202];
endrule
rule s1204(sum_count == 1204);
  total_sum <= total_sum + cache[1203];
endrule
rule s1205(sum_count == 1205);
  total_sum <= total_sum + cache[1204];
endrule
rule s1206(sum_count == 1206);
  total_sum <= total_sum + cache[1205];
endrule
rule s1207(sum_count == 1207);
  total_sum <= total_sum + cache[1206];
endrule
rule s1208(sum_count == 1208);
  total_sum <= total_sum + cache[1207];
endrule
rule s1209(sum_count == 1209);
  total_sum <= total_sum + cache[1208];
endrule
rule s1210(sum_count == 1210);
  total_sum <= total_sum + cache[1209];
endrule
rule s1211(sum_count == 1211);
  total_sum <= total_sum + cache[1210];
endrule
rule s1212(sum_count == 1212);
  total_sum <= total_sum + cache[1211];
endrule
rule s1213(sum_count == 1213);
  total_sum <= total_sum + cache[1212];
endrule
rule s1214(sum_count == 1214);
  total_sum <= total_sum + cache[1213];
endrule
rule s1215(sum_count == 1215);
  total_sum <= total_sum + cache[1214];
endrule
rule s1216(sum_count == 1216);
  total_sum <= total_sum + cache[1215];
endrule
rule s1217(sum_count == 1217);
  total_sum <= total_sum + cache[1216];
endrule
rule s1218(sum_count == 1218);
  total_sum <= total_sum + cache[1217];
endrule
rule s1219(sum_count == 1219);
  total_sum <= total_sum + cache[1218];
endrule
rule s1220(sum_count == 1220);
  total_sum <= total_sum + cache[1219];
endrule
rule s1221(sum_count == 1221);
  total_sum <= total_sum + cache[1220];
endrule
rule s1222(sum_count == 1222);
  total_sum <= total_sum + cache[1221];
endrule
rule s1223(sum_count == 1223);
  total_sum <= total_sum + cache[1222];
endrule
rule s1224(sum_count == 1224);
  total_sum <= total_sum + cache[1223];
endrule
rule s1225(sum_count == 1225);
  total_sum <= total_sum + cache[1224];
endrule
rule s1226(sum_count == 1226);
  total_sum <= total_sum + cache[1225];
endrule
rule s1227(sum_count == 1227);
  total_sum <= total_sum + cache[1226];
endrule
rule s1228(sum_count == 1228);
  total_sum <= total_sum + cache[1227];
endrule
rule s1229(sum_count == 1229);
  total_sum <= total_sum + cache[1228];
endrule
rule s1230(sum_count == 1230);
  total_sum <= total_sum + cache[1229];
endrule
rule s1231(sum_count == 1231);
  total_sum <= total_sum + cache[1230];
endrule
rule s1232(sum_count == 1232);
  total_sum <= total_sum + cache[1231];
endrule
rule s1233(sum_count == 1233);
  total_sum <= total_sum + cache[1232];
endrule
rule s1234(sum_count == 1234);
  total_sum <= total_sum + cache[1233];
endrule
rule s1235(sum_count == 1235);
  total_sum <= total_sum + cache[1234];
endrule
rule s1236(sum_count == 1236);
  total_sum <= total_sum + cache[1235];
endrule
rule s1237(sum_count == 1237);
  total_sum <= total_sum + cache[1236];
endrule
rule s1238(sum_count == 1238);
  total_sum <= total_sum + cache[1237];
endrule
rule s1239(sum_count == 1239);
  total_sum <= total_sum + cache[1238];
endrule
rule s1240(sum_count == 1240);
  total_sum <= total_sum + cache[1239];
endrule
rule s1241(sum_count == 1241);
  total_sum <= total_sum + cache[1240];
endrule
rule s1242(sum_count == 1242);
  total_sum <= total_sum + cache[1241];
endrule
rule s1243(sum_count == 1243);
  total_sum <= total_sum + cache[1242];
endrule
rule s1244(sum_count == 1244);
  total_sum <= total_sum + cache[1243];
endrule
rule s1245(sum_count == 1245);
  total_sum <= total_sum + cache[1244];
endrule
rule s1246(sum_count == 1246);
  total_sum <= total_sum + cache[1245];
endrule
rule s1247(sum_count == 1247);
  total_sum <= total_sum + cache[1246];
endrule
rule s1248(sum_count == 1248);
  total_sum <= total_sum + cache[1247];
endrule
rule s1249(sum_count == 1249);
  total_sum <= total_sum + cache[1248];
endrule
rule s1250(sum_count == 1250);
  total_sum <= total_sum + cache[1249];
endrule
rule s1251(sum_count == 1251);
  total_sum <= total_sum + cache[1250];
endrule
rule s1252(sum_count == 1252);
  total_sum <= total_sum + cache[1251];
endrule
rule s1253(sum_count == 1253);
  total_sum <= total_sum + cache[1252];
endrule
rule s1254(sum_count == 1254);
  total_sum <= total_sum + cache[1253];
endrule
rule s1255(sum_count == 1255);
  total_sum <= total_sum + cache[1254];
endrule
rule s1256(sum_count == 1256);
  total_sum <= total_sum + cache[1255];
endrule
rule s1257(sum_count == 1257);
  total_sum <= total_sum + cache[1256];
endrule
rule s1258(sum_count == 1258);
  total_sum <= total_sum + cache[1257];
endrule
rule s1259(sum_count == 1259);
  total_sum <= total_sum + cache[1258];
endrule
rule s1260(sum_count == 1260);
  total_sum <= total_sum + cache[1259];
endrule
rule s1261(sum_count == 1261);
  total_sum <= total_sum + cache[1260];
endrule
rule s1262(sum_count == 1262);
  total_sum <= total_sum + cache[1261];
endrule
rule s1263(sum_count == 1263);
  total_sum <= total_sum + cache[1262];
endrule
rule s1264(sum_count == 1264);
  total_sum <= total_sum + cache[1263];
endrule
rule s1265(sum_count == 1265);
  total_sum <= total_sum + cache[1264];
endrule
rule s1266(sum_count == 1266);
  total_sum <= total_sum + cache[1265];
endrule
rule s1267(sum_count == 1267);
  total_sum <= total_sum + cache[1266];
endrule
rule s1268(sum_count == 1268);
  total_sum <= total_sum + cache[1267];
endrule
rule s1269(sum_count == 1269);
  total_sum <= total_sum + cache[1268];
endrule
rule s1270(sum_count == 1270);
  total_sum <= total_sum + cache[1269];
endrule
rule s1271(sum_count == 1271);
  total_sum <= total_sum + cache[1270];
endrule
rule s1272(sum_count == 1272);
  total_sum <= total_sum + cache[1271];
endrule
rule s1273(sum_count == 1273);
  total_sum <= total_sum + cache[1272];
endrule
rule s1274(sum_count == 1274);
  total_sum <= total_sum + cache[1273];
endrule
rule s1275(sum_count == 1275);
  total_sum <= total_sum + cache[1274];
endrule
rule s1276(sum_count == 1276);
  total_sum <= total_sum + cache[1275];
endrule
rule s1277(sum_count == 1277);
  total_sum <= total_sum + cache[1276];
endrule
rule s1278(sum_count == 1278);
  total_sum <= total_sum + cache[1277];
endrule
rule s1279(sum_count == 1279);
  total_sum <= total_sum + cache[1278];
endrule
rule s1280(sum_count == 1280);
  total_sum <= total_sum + cache[1279];
endrule
rule s1281(sum_count == 1281);
  total_sum <= total_sum + cache[1280];
endrule
rule s1282(sum_count == 1282);
  total_sum <= total_sum + cache[1281];
endrule
rule s1283(sum_count == 1283);
  total_sum <= total_sum + cache[1282];
endrule
rule s1284(sum_count == 1284);
  total_sum <= total_sum + cache[1283];
endrule
rule s1285(sum_count == 1285);
  total_sum <= total_sum + cache[1284];
endrule
rule s1286(sum_count == 1286);
  total_sum <= total_sum + cache[1285];
endrule
rule s1287(sum_count == 1287);
  total_sum <= total_sum + cache[1286];
endrule
rule s1288(sum_count == 1288);
  total_sum <= total_sum + cache[1287];
endrule
rule s1289(sum_count == 1289);
  total_sum <= total_sum + cache[1288];
endrule
rule s1290(sum_count == 1290);
  total_sum <= total_sum + cache[1289];
endrule
rule s1291(sum_count == 1291);
  total_sum <= total_sum + cache[1290];
endrule
rule s1292(sum_count == 1292);
  total_sum <= total_sum + cache[1291];
endrule
rule s1293(sum_count == 1293);
  total_sum <= total_sum + cache[1292];
endrule
rule s1294(sum_count == 1294);
  total_sum <= total_sum + cache[1293];
endrule
rule s1295(sum_count == 1295);
  total_sum <= total_sum + cache[1294];
endrule
rule s1296(sum_count == 1296);
  total_sum <= total_sum + cache[1295];
endrule
rule s1297(sum_count == 1297);
  total_sum <= total_sum + cache[1296];
endrule
rule s1298(sum_count == 1298);
  total_sum <= total_sum + cache[1297];
endrule
rule s1299(sum_count == 1299);
  total_sum <= total_sum + cache[1298];
endrule
rule s1300(sum_count == 1300);
  total_sum <= total_sum + cache[1299];
endrule
rule s1301(sum_count == 1301);
  total_sum <= total_sum + cache[1300];
endrule
rule s1302(sum_count == 1302);
  total_sum <= total_sum + cache[1301];
endrule
rule s1303(sum_count == 1303);
  total_sum <= total_sum + cache[1302];
endrule
rule s1304(sum_count == 1304);
  total_sum <= total_sum + cache[1303];
endrule
rule s1305(sum_count == 1305);
  total_sum <= total_sum + cache[1304];
endrule
rule s1306(sum_count == 1306);
  total_sum <= total_sum + cache[1305];
endrule
rule s1307(sum_count == 1307);
  total_sum <= total_sum + cache[1306];
endrule
rule s1308(sum_count == 1308);
  total_sum <= total_sum + cache[1307];
endrule
rule s1309(sum_count == 1309);
  total_sum <= total_sum + cache[1308];
endrule
rule s1310(sum_count == 1310);
  total_sum <= total_sum + cache[1309];
endrule
rule s1311(sum_count == 1311);
  total_sum <= total_sum + cache[1310];
endrule
rule s1312(sum_count == 1312);
  total_sum <= total_sum + cache[1311];
endrule
rule s1313(sum_count == 1313);
  total_sum <= total_sum + cache[1312];
endrule
rule s1314(sum_count == 1314);
  total_sum <= total_sum + cache[1313];
endrule
rule s1315(sum_count == 1315);
  total_sum <= total_sum + cache[1314];
endrule
rule s1316(sum_count == 1316);
  total_sum <= total_sum + cache[1315];
endrule
rule s1317(sum_count == 1317);
  total_sum <= total_sum + cache[1316];
endrule
rule s1318(sum_count == 1318);
  total_sum <= total_sum + cache[1317];
endrule
rule s1319(sum_count == 1319);
  total_sum <= total_sum + cache[1318];
endrule
rule s1320(sum_count == 1320);
  total_sum <= total_sum + cache[1319];
endrule
rule s1321(sum_count == 1321);
  total_sum <= total_sum + cache[1320];
endrule
rule s1322(sum_count == 1322);
  total_sum <= total_sum + cache[1321];
endrule
rule s1323(sum_count == 1323);
  total_sum <= total_sum + cache[1322];
endrule
rule s1324(sum_count == 1324);
  total_sum <= total_sum + cache[1323];
endrule
rule s1325(sum_count == 1325);
  total_sum <= total_sum + cache[1324];
endrule
rule s1326(sum_count == 1326);
  total_sum <= total_sum + cache[1325];
endrule
rule s1327(sum_count == 1327);
  total_sum <= total_sum + cache[1326];
endrule
rule s1328(sum_count == 1328);
  total_sum <= total_sum + cache[1327];
endrule
rule s1329(sum_count == 1329);
  total_sum <= total_sum + cache[1328];
endrule
rule s1330(sum_count == 1330);
  total_sum <= total_sum + cache[1329];
endrule
rule s1331(sum_count == 1331);
  total_sum <= total_sum + cache[1330];
endrule
rule s1332(sum_count == 1332);
  total_sum <= total_sum + cache[1331];
endrule
rule s1333(sum_count == 1333);
  total_sum <= total_sum + cache[1332];
endrule
rule s1334(sum_count == 1334);
  total_sum <= total_sum + cache[1333];
endrule
rule s1335(sum_count == 1335);
  total_sum <= total_sum + cache[1334];
endrule
rule s1336(sum_count == 1336);
  total_sum <= total_sum + cache[1335];
endrule
rule s1337(sum_count == 1337);
  total_sum <= total_sum + cache[1336];
endrule
rule s1338(sum_count == 1338);
  total_sum <= total_sum + cache[1337];
endrule
rule s1339(sum_count == 1339);
  total_sum <= total_sum + cache[1338];
endrule
rule s1340(sum_count == 1340);
  total_sum <= total_sum + cache[1339];
endrule
rule s1341(sum_count == 1341);
  total_sum <= total_sum + cache[1340];
endrule
rule s1342(sum_count == 1342);
  total_sum <= total_sum + cache[1341];
endrule
rule s1343(sum_count == 1343);
  total_sum <= total_sum + cache[1342];
endrule
rule s1344(sum_count == 1344);
  total_sum <= total_sum + cache[1343];
endrule
rule s1345(sum_count == 1345);
  total_sum <= total_sum + cache[1344];
endrule
rule s1346(sum_count == 1346);
  total_sum <= total_sum + cache[1345];
endrule
rule s1347(sum_count == 1347);
  total_sum <= total_sum + cache[1346];
endrule
rule s1348(sum_count == 1348);
  total_sum <= total_sum + cache[1347];
endrule
rule s1349(sum_count == 1349);
  total_sum <= total_sum + cache[1348];
endrule
rule s1350(sum_count == 1350);
  total_sum <= total_sum + cache[1349];
endrule
rule s1351(sum_count == 1351);
  total_sum <= total_sum + cache[1350];
endrule
rule s1352(sum_count == 1352);
  total_sum <= total_sum + cache[1351];
endrule
rule s1353(sum_count == 1353);
  total_sum <= total_sum + cache[1352];
endrule
rule s1354(sum_count == 1354);
  total_sum <= total_sum + cache[1353];
endrule
rule s1355(sum_count == 1355);
  total_sum <= total_sum + cache[1354];
endrule
rule s1356(sum_count == 1356);
  total_sum <= total_sum + cache[1355];
endrule
rule s1357(sum_count == 1357);
  total_sum <= total_sum + cache[1356];
endrule
rule s1358(sum_count == 1358);
  total_sum <= total_sum + cache[1357];
endrule
rule s1359(sum_count == 1359);
  total_sum <= total_sum + cache[1358];
endrule
rule s1360(sum_count == 1360);
  total_sum <= total_sum + cache[1359];
endrule
rule s1361(sum_count == 1361);
  total_sum <= total_sum + cache[1360];
endrule
rule s1362(sum_count == 1362);
  total_sum <= total_sum + cache[1361];
endrule
rule s1363(sum_count == 1363);
  total_sum <= total_sum + cache[1362];
endrule
rule s1364(sum_count == 1364);
  total_sum <= total_sum + cache[1363];
endrule
rule s1365(sum_count == 1365);
  total_sum <= total_sum + cache[1364];
endrule
rule s1366(sum_count == 1366);
  total_sum <= total_sum + cache[1365];
endrule
rule s1367(sum_count == 1367);
  total_sum <= total_sum + cache[1366];
endrule
rule s1368(sum_count == 1368);
  total_sum <= total_sum + cache[1367];
endrule
rule s1369(sum_count == 1369);
  total_sum <= total_sum + cache[1368];
endrule
rule s1370(sum_count == 1370);
  total_sum <= total_sum + cache[1369];
endrule
rule s1371(sum_count == 1371);
  total_sum <= total_sum + cache[1370];
endrule
rule s1372(sum_count == 1372);
  total_sum <= total_sum + cache[1371];
endrule
rule s1373(sum_count == 1373);
  total_sum <= total_sum + cache[1372];
endrule
rule s1374(sum_count == 1374);
  total_sum <= total_sum + cache[1373];
endrule
rule s1375(sum_count == 1375);
  total_sum <= total_sum + cache[1374];
endrule
rule s1376(sum_count == 1376);
  total_sum <= total_sum + cache[1375];
endrule
rule s1377(sum_count == 1377);
  total_sum <= total_sum + cache[1376];
endrule
rule s1378(sum_count == 1378);
  total_sum <= total_sum + cache[1377];
endrule
rule s1379(sum_count == 1379);
  total_sum <= total_sum + cache[1378];
endrule
rule s1380(sum_count == 1380);
  total_sum <= total_sum + cache[1379];
endrule
rule s1381(sum_count == 1381);
  total_sum <= total_sum + cache[1380];
endrule
rule s1382(sum_count == 1382);
  total_sum <= total_sum + cache[1381];
endrule
rule s1383(sum_count == 1383);
  total_sum <= total_sum + cache[1382];
endrule
rule s1384(sum_count == 1384);
  total_sum <= total_sum + cache[1383];
endrule
rule s1385(sum_count == 1385);
  total_sum <= total_sum + cache[1384];
endrule
rule s1386(sum_count == 1386);
  total_sum <= total_sum + cache[1385];
endrule
rule s1387(sum_count == 1387);
  total_sum <= total_sum + cache[1386];
endrule
rule s1388(sum_count == 1388);
  total_sum <= total_sum + cache[1387];
endrule
rule s1389(sum_count == 1389);
  total_sum <= total_sum + cache[1388];
endrule
rule s1390(sum_count == 1390);
  total_sum <= total_sum + cache[1389];
endrule
rule s1391(sum_count == 1391);
  total_sum <= total_sum + cache[1390];
endrule
rule s1392(sum_count == 1392);
  total_sum <= total_sum + cache[1391];
endrule
rule s1393(sum_count == 1393);
  total_sum <= total_sum + cache[1392];
endrule
rule s1394(sum_count == 1394);
  total_sum <= total_sum + cache[1393];
endrule
rule s1395(sum_count == 1395);
  total_sum <= total_sum + cache[1394];
endrule
rule s1396(sum_count == 1396);
  total_sum <= total_sum + cache[1395];
endrule
rule s1397(sum_count == 1397);
  total_sum <= total_sum + cache[1396];
endrule
rule s1398(sum_count == 1398);
  total_sum <= total_sum + cache[1397];
endrule
rule s1399(sum_count == 1399);
  total_sum <= total_sum + cache[1398];
endrule
rule s1400(sum_count == 1400);
  total_sum <= total_sum + cache[1399];
endrule
rule s1401(sum_count == 1401);
  total_sum <= total_sum + cache[1400];
endrule
rule s1402(sum_count == 1402);
  total_sum <= total_sum + cache[1401];
endrule
rule s1403(sum_count == 1403);
  total_sum <= total_sum + cache[1402];
endrule
rule s1404(sum_count == 1404);
  total_sum <= total_sum + cache[1403];
endrule
rule s1405(sum_count == 1405);
  total_sum <= total_sum + cache[1404];
endrule
rule s1406(sum_count == 1406);
  total_sum <= total_sum + cache[1405];
endrule
rule s1407(sum_count == 1407);
  total_sum <= total_sum + cache[1406];
endrule
rule s1408(sum_count == 1408);
  total_sum <= total_sum + cache[1407];
endrule
rule s1409(sum_count == 1409);
  total_sum <= total_sum + cache[1408];
endrule
rule s1410(sum_count == 1410);
  total_sum <= total_sum + cache[1409];
endrule
rule s1411(sum_count == 1411);
  total_sum <= total_sum + cache[1410];
endrule
rule s1412(sum_count == 1412);
  total_sum <= total_sum + cache[1411];
endrule
rule s1413(sum_count == 1413);
  total_sum <= total_sum + cache[1412];
endrule
rule s1414(sum_count == 1414);
  total_sum <= total_sum + cache[1413];
endrule
rule s1415(sum_count == 1415);
  total_sum <= total_sum + cache[1414];
endrule
rule s1416(sum_count == 1416);
  total_sum <= total_sum + cache[1415];
endrule
rule s1417(sum_count == 1417);
  total_sum <= total_sum + cache[1416];
endrule
rule s1418(sum_count == 1418);
  total_sum <= total_sum + cache[1417];
endrule
rule s1419(sum_count == 1419);
  total_sum <= total_sum + cache[1418];
endrule
rule s1420(sum_count == 1420);
  total_sum <= total_sum + cache[1419];
endrule
rule s1421(sum_count == 1421);
  total_sum <= total_sum + cache[1420];
endrule
rule s1422(sum_count == 1422);
  total_sum <= total_sum + cache[1421];
endrule
rule s1423(sum_count == 1423);
  total_sum <= total_sum + cache[1422];
endrule
rule s1424(sum_count == 1424);
  total_sum <= total_sum + cache[1423];
endrule
rule s1425(sum_count == 1425);
  total_sum <= total_sum + cache[1424];
endrule
rule s1426(sum_count == 1426);
  total_sum <= total_sum + cache[1425];
endrule
rule s1427(sum_count == 1427);
  total_sum <= total_sum + cache[1426];
endrule
rule s1428(sum_count == 1428);
  total_sum <= total_sum + cache[1427];
endrule
rule s1429(sum_count == 1429);
  total_sum <= total_sum + cache[1428];
endrule
rule s1430(sum_count == 1430);
  total_sum <= total_sum + cache[1429];
endrule
rule s1431(sum_count == 1431);
  total_sum <= total_sum + cache[1430];
endrule
rule s1432(sum_count == 1432);
  total_sum <= total_sum + cache[1431];
endrule
rule s1433(sum_count == 1433);
  total_sum <= total_sum + cache[1432];
endrule
rule s1434(sum_count == 1434);
  total_sum <= total_sum + cache[1433];
endrule
rule s1435(sum_count == 1435);
  total_sum <= total_sum + cache[1434];
endrule
rule s1436(sum_count == 1436);
  total_sum <= total_sum + cache[1435];
endrule
rule s1437(sum_count == 1437);
  total_sum <= total_sum + cache[1436];
endrule
rule s1438(sum_count == 1438);
  total_sum <= total_sum + cache[1437];
endrule
rule s1439(sum_count == 1439);
  total_sum <= total_sum + cache[1438];
endrule
rule s1440(sum_count == 1440);
  total_sum <= total_sum + cache[1439];
endrule
rule s1441(sum_count == 1441);
  total_sum <= total_sum + cache[1440];
endrule
rule s1442(sum_count == 1442);
  total_sum <= total_sum + cache[1441];
endrule
rule s1443(sum_count == 1443);
  total_sum <= total_sum + cache[1442];
endrule
rule s1444(sum_count == 1444);
  total_sum <= total_sum + cache[1443];
endrule
rule s1445(sum_count == 1445);
  total_sum <= total_sum + cache[1444];
endrule
rule s1446(sum_count == 1446);
  total_sum <= total_sum + cache[1445];
endrule
rule s1447(sum_count == 1447);
  total_sum <= total_sum + cache[1446];
endrule
rule s1448(sum_count == 1448);
  total_sum <= total_sum + cache[1447];
endrule
rule s1449(sum_count == 1449);
  total_sum <= total_sum + cache[1448];
endrule
rule s1450(sum_count == 1450);
  total_sum <= total_sum + cache[1449];
endrule
rule s1451(sum_count == 1451);
  total_sum <= total_sum + cache[1450];
endrule
rule s1452(sum_count == 1452);
  total_sum <= total_sum + cache[1451];
endrule
rule s1453(sum_count == 1453);
  total_sum <= total_sum + cache[1452];
endrule
rule s1454(sum_count == 1454);
  total_sum <= total_sum + cache[1453];
endrule
rule s1455(sum_count == 1455);
  total_sum <= total_sum + cache[1454];
endrule
rule s1456(sum_count == 1456);
  total_sum <= total_sum + cache[1455];
endrule
rule s1457(sum_count == 1457);
  total_sum <= total_sum + cache[1456];
endrule
rule s1458(sum_count == 1458);
  total_sum <= total_sum + cache[1457];
endrule
rule s1459(sum_count == 1459);
  total_sum <= total_sum + cache[1458];
endrule
rule s1460(sum_count == 1460);
  total_sum <= total_sum + cache[1459];
endrule
rule s1461(sum_count == 1461);
  total_sum <= total_sum + cache[1460];
endrule
rule s1462(sum_count == 1462);
  total_sum <= total_sum + cache[1461];
endrule
rule s1463(sum_count == 1463);
  total_sum <= total_sum + cache[1462];
endrule
rule s1464(sum_count == 1464);
  total_sum <= total_sum + cache[1463];
endrule
rule s1465(sum_count == 1465);
  total_sum <= total_sum + cache[1464];
endrule
rule s1466(sum_count == 1466);
  total_sum <= total_sum + cache[1465];
endrule
rule s1467(sum_count == 1467);
  total_sum <= total_sum + cache[1466];
endrule
rule s1468(sum_count == 1468);
  total_sum <= total_sum + cache[1467];
endrule
rule s1469(sum_count == 1469);
  total_sum <= total_sum + cache[1468];
endrule
rule s1470(sum_count == 1470);
  total_sum <= total_sum + cache[1469];
endrule
rule s1471(sum_count == 1471);
  total_sum <= total_sum + cache[1470];
endrule
rule s1472(sum_count == 1472);
  total_sum <= total_sum + cache[1471];
endrule
rule s1473(sum_count == 1473);
  total_sum <= total_sum + cache[1472];
endrule
rule s1474(sum_count == 1474);
  total_sum <= total_sum + cache[1473];
endrule
rule s1475(sum_count == 1475);
  total_sum <= total_sum + cache[1474];
endrule
rule s1476(sum_count == 1476);
  total_sum <= total_sum + cache[1475];
endrule
rule s1477(sum_count == 1477);
  total_sum <= total_sum + cache[1476];
endrule
rule s1478(sum_count == 1478);
  total_sum <= total_sum + cache[1477];
endrule
rule s1479(sum_count == 1479);
  total_sum <= total_sum + cache[1478];
endrule
rule s1480(sum_count == 1480);
  total_sum <= total_sum + cache[1479];
endrule
rule s1481(sum_count == 1481);
  total_sum <= total_sum + cache[1480];
endrule
rule s1482(sum_count == 1482);
  total_sum <= total_sum + cache[1481];
endrule
rule s1483(sum_count == 1483);
  total_sum <= total_sum + cache[1482];
endrule
rule s1484(sum_count == 1484);
  total_sum <= total_sum + cache[1483];
endrule
rule s1485(sum_count == 1485);
  total_sum <= total_sum + cache[1484];
endrule
rule s1486(sum_count == 1486);
  total_sum <= total_sum + cache[1485];
endrule
rule s1487(sum_count == 1487);
  total_sum <= total_sum + cache[1486];
endrule
rule s1488(sum_count == 1488);
  total_sum <= total_sum + cache[1487];
endrule
rule s1489(sum_count == 1489);
  total_sum <= total_sum + cache[1488];
endrule
rule s1490(sum_count == 1490);
  total_sum <= total_sum + cache[1489];
endrule
rule s1491(sum_count == 1491);
  total_sum <= total_sum + cache[1490];
endrule
rule s1492(sum_count == 1492);
  total_sum <= total_sum + cache[1491];
endrule
rule s1493(sum_count == 1493);
  total_sum <= total_sum + cache[1492];
endrule
rule s1494(sum_count == 1494);
  total_sum <= total_sum + cache[1493];
endrule
rule s1495(sum_count == 1495);
  total_sum <= total_sum + cache[1494];
endrule
rule s1496(sum_count == 1496);
  total_sum <= total_sum + cache[1495];
endrule
rule s1497(sum_count == 1497);
  total_sum <= total_sum + cache[1496];
endrule
rule s1498(sum_count == 1498);
  total_sum <= total_sum + cache[1497];
endrule
rule s1499(sum_count == 1499);
  total_sum <= total_sum + cache[1498];
endrule
rule s1500(sum_count == 1500);
  total_sum <= total_sum + cache[1499];
endrule
rule s1501(sum_count == 1501);
  total_sum <= total_sum + cache[1500];
endrule
rule s1502(sum_count == 1502);
  total_sum <= total_sum + cache[1501];
endrule
rule s1503(sum_count == 1503);
  total_sum <= total_sum + cache[1502];
endrule
rule s1504(sum_count == 1504);
  total_sum <= total_sum + cache[1503];
endrule
rule s1505(sum_count == 1505);
  total_sum <= total_sum + cache[1504];
endrule
rule s1506(sum_count == 1506);
  total_sum <= total_sum + cache[1505];
endrule
rule s1507(sum_count == 1507);
  total_sum <= total_sum + cache[1506];
endrule
rule s1508(sum_count == 1508);
  total_sum <= total_sum + cache[1507];
endrule
rule s1509(sum_count == 1509);
  total_sum <= total_sum + cache[1508];
endrule
rule s1510(sum_count == 1510);
  total_sum <= total_sum + cache[1509];
endrule
rule s1511(sum_count == 1511);
  total_sum <= total_sum + cache[1510];
endrule
rule s1512(sum_count == 1512);
  total_sum <= total_sum + cache[1511];
endrule
rule s1513(sum_count == 1513);
  total_sum <= total_sum + cache[1512];
endrule
rule s1514(sum_count == 1514);
  total_sum <= total_sum + cache[1513];
endrule
rule s1515(sum_count == 1515);
  total_sum <= total_sum + cache[1514];
endrule
rule s1516(sum_count == 1516);
  total_sum <= total_sum + cache[1515];
endrule
rule s1517(sum_count == 1517);
  total_sum <= total_sum + cache[1516];
endrule
rule s1518(sum_count == 1518);
  total_sum <= total_sum + cache[1517];
endrule
rule s1519(sum_count == 1519);
  total_sum <= total_sum + cache[1518];
endrule
rule s1520(sum_count == 1520);
  total_sum <= total_sum + cache[1519];
endrule
rule s1521(sum_count == 1521);
  total_sum <= total_sum + cache[1520];
endrule
rule s1522(sum_count == 1522);
  total_sum <= total_sum + cache[1521];
endrule
rule s1523(sum_count == 1523);
  total_sum <= total_sum + cache[1522];
endrule
rule s1524(sum_count == 1524);
  total_sum <= total_sum + cache[1523];
endrule
rule s1525(sum_count == 1525);
  total_sum <= total_sum + cache[1524];
endrule
rule s1526(sum_count == 1526);
  total_sum <= total_sum + cache[1525];
endrule
rule s1527(sum_count == 1527);
  total_sum <= total_sum + cache[1526];
endrule
rule s1528(sum_count == 1528);
  total_sum <= total_sum + cache[1527];
endrule
rule s1529(sum_count == 1529);
  total_sum <= total_sum + cache[1528];
endrule
rule s1530(sum_count == 1530);
  total_sum <= total_sum + cache[1529];
endrule
rule s1531(sum_count == 1531);
  total_sum <= total_sum + cache[1530];
endrule
rule s1532(sum_count == 1532);
  total_sum <= total_sum + cache[1531];
endrule
rule s1533(sum_count == 1533);
  total_sum <= total_sum + cache[1532];
endrule
rule s1534(sum_count == 1534);
  total_sum <= total_sum + cache[1533];
endrule
rule s1535(sum_count == 1535);
  total_sum <= total_sum + cache[1534];
endrule
rule s1536(sum_count == 1536);
  total_sum <= total_sum + cache[1535];
endrule
rule s1537(sum_count == 1537);
  total_sum <= total_sum + cache[1536];
endrule
rule s1538(sum_count == 1538);
  total_sum <= total_sum + cache[1537];
endrule
rule s1539(sum_count == 1539);
  total_sum <= total_sum + cache[1538];
endrule
rule s1540(sum_count == 1540);
  total_sum <= total_sum + cache[1539];
endrule
rule s1541(sum_count == 1541);
  total_sum <= total_sum + cache[1540];
endrule
rule s1542(sum_count == 1542);
  total_sum <= total_sum + cache[1541];
endrule
rule s1543(sum_count == 1543);
  total_sum <= total_sum + cache[1542];
endrule
rule s1544(sum_count == 1544);
  total_sum <= total_sum + cache[1543];
endrule
rule s1545(sum_count == 1545);
  total_sum <= total_sum + cache[1544];
endrule
rule s1546(sum_count == 1546);
  total_sum <= total_sum + cache[1545];
endrule
rule s1547(sum_count == 1547);
  total_sum <= total_sum + cache[1546];
endrule
rule s1548(sum_count == 1548);
  total_sum <= total_sum + cache[1547];
endrule
rule s1549(sum_count == 1549);
  total_sum <= total_sum + cache[1548];
endrule
rule s1550(sum_count == 1550);
  total_sum <= total_sum + cache[1549];
endrule
rule s1551(sum_count == 1551);
  total_sum <= total_sum + cache[1550];
endrule
rule s1552(sum_count == 1552);
  total_sum <= total_sum + cache[1551];
endrule
rule s1553(sum_count == 1553);
  total_sum <= total_sum + cache[1552];
endrule
rule s1554(sum_count == 1554);
  total_sum <= total_sum + cache[1553];
endrule
rule s1555(sum_count == 1555);
  total_sum <= total_sum + cache[1554];
endrule
rule s1556(sum_count == 1556);
  total_sum <= total_sum + cache[1555];
endrule
rule s1557(sum_count == 1557);
  total_sum <= total_sum + cache[1556];
endrule
rule s1558(sum_count == 1558);
  total_sum <= total_sum + cache[1557];
endrule
rule s1559(sum_count == 1559);
  total_sum <= total_sum + cache[1558];
endrule
rule s1560(sum_count == 1560);
  total_sum <= total_sum + cache[1559];
endrule
rule s1561(sum_count == 1561);
  total_sum <= total_sum + cache[1560];
endrule
rule s1562(sum_count == 1562);
  total_sum <= total_sum + cache[1561];
endrule
rule s1563(sum_count == 1563);
  total_sum <= total_sum + cache[1562];
endrule
rule s1564(sum_count == 1564);
  total_sum <= total_sum + cache[1563];
endrule
rule s1565(sum_count == 1565);
  total_sum <= total_sum + cache[1564];
endrule
rule s1566(sum_count == 1566);
  total_sum <= total_sum + cache[1565];
endrule
rule s1567(sum_count == 1567);
  total_sum <= total_sum + cache[1566];
endrule
rule s1568(sum_count == 1568);
  total_sum <= total_sum + cache[1567];
endrule
rule s1569(sum_count == 1569);
  total_sum <= total_sum + cache[1568];
endrule
rule s1570(sum_count == 1570);
  total_sum <= total_sum + cache[1569];
endrule
rule s1571(sum_count == 1571);
  total_sum <= total_sum + cache[1570];
endrule
rule s1572(sum_count == 1572);
  total_sum <= total_sum + cache[1571];
endrule
rule s1573(sum_count == 1573);
  total_sum <= total_sum + cache[1572];
endrule
rule s1574(sum_count == 1574);
  total_sum <= total_sum + cache[1573];
endrule
rule s1575(sum_count == 1575);
  total_sum <= total_sum + cache[1574];
endrule
rule s1576(sum_count == 1576);
  total_sum <= total_sum + cache[1575];
endrule
rule s1577(sum_count == 1577);
  total_sum <= total_sum + cache[1576];
endrule
rule s1578(sum_count == 1578);
  total_sum <= total_sum + cache[1577];
endrule
rule s1579(sum_count == 1579);
  total_sum <= total_sum + cache[1578];
endrule
rule s1580(sum_count == 1580);
  total_sum <= total_sum + cache[1579];
endrule
rule s1581(sum_count == 1581);
  total_sum <= total_sum + cache[1580];
endrule
rule s1582(sum_count == 1582);
  total_sum <= total_sum + cache[1581];
endrule
rule s1583(sum_count == 1583);
  total_sum <= total_sum + cache[1582];
endrule
rule s1584(sum_count == 1584);
  total_sum <= total_sum + cache[1583];
endrule
rule s1585(sum_count == 1585);
  total_sum <= total_sum + cache[1584];
endrule
rule s1586(sum_count == 1586);
  total_sum <= total_sum + cache[1585];
endrule
rule s1587(sum_count == 1587);
  total_sum <= total_sum + cache[1586];
endrule
rule s1588(sum_count == 1588);
  total_sum <= total_sum + cache[1587];
endrule
rule s1589(sum_count == 1589);
  total_sum <= total_sum + cache[1588];
endrule
rule s1590(sum_count == 1590);
  total_sum <= total_sum + cache[1589];
endrule
rule s1591(sum_count == 1591);
  total_sum <= total_sum + cache[1590];
endrule
rule s1592(sum_count == 1592);
  total_sum <= total_sum + cache[1591];
endrule
rule s1593(sum_count == 1593);
  total_sum <= total_sum + cache[1592];
endrule
rule s1594(sum_count == 1594);
  total_sum <= total_sum + cache[1593];
endrule
rule s1595(sum_count == 1595);
  total_sum <= total_sum + cache[1594];
endrule
rule s1596(sum_count == 1596);
  total_sum <= total_sum + cache[1595];
endrule
rule s1597(sum_count == 1597);
  total_sum <= total_sum + cache[1596];
endrule
rule s1598(sum_count == 1598);
  total_sum <= total_sum + cache[1597];
endrule
rule s1599(sum_count == 1599);
  total_sum <= total_sum + cache[1598];
endrule
rule s1600(sum_count == 1600);
  total_sum <= total_sum + cache[1599];
endrule
rule s1601(sum_count == 1601);
  total_sum <= total_sum + cache[1600];
endrule
rule s1602(sum_count == 1602);
  total_sum <= total_sum + cache[1601];
endrule
rule s1603(sum_count == 1603);
  total_sum <= total_sum + cache[1602];
endrule
rule s1604(sum_count == 1604);
  total_sum <= total_sum + cache[1603];
endrule
rule s1605(sum_count == 1605);
  total_sum <= total_sum + cache[1604];
endrule
rule s1606(sum_count == 1606);
  total_sum <= total_sum + cache[1605];
endrule
rule s1607(sum_count == 1607);
  total_sum <= total_sum + cache[1606];
endrule
rule s1608(sum_count == 1608);
  total_sum <= total_sum + cache[1607];
endrule
rule s1609(sum_count == 1609);
  total_sum <= total_sum + cache[1608];
endrule
rule s1610(sum_count == 1610);
  total_sum <= total_sum + cache[1609];
endrule
rule s1611(sum_count == 1611);
  total_sum <= total_sum + cache[1610];
endrule
rule s1612(sum_count == 1612);
  total_sum <= total_sum + cache[1611];
endrule
rule s1613(sum_count == 1613);
  total_sum <= total_sum + cache[1612];
endrule
rule s1614(sum_count == 1614);
  total_sum <= total_sum + cache[1613];
endrule
rule s1615(sum_count == 1615);
  total_sum <= total_sum + cache[1614];
endrule
rule s1616(sum_count == 1616);
  total_sum <= total_sum + cache[1615];
endrule
rule s1617(sum_count == 1617);
  total_sum <= total_sum + cache[1616];
endrule
rule s1618(sum_count == 1618);
  total_sum <= total_sum + cache[1617];
endrule
rule s1619(sum_count == 1619);
  total_sum <= total_sum + cache[1618];
endrule
rule s1620(sum_count == 1620);
  total_sum <= total_sum + cache[1619];
endrule
rule s1621(sum_count == 1621);
  total_sum <= total_sum + cache[1620];
endrule
rule s1622(sum_count == 1622);
  total_sum <= total_sum + cache[1621];
endrule
rule s1623(sum_count == 1623);
  total_sum <= total_sum + cache[1622];
endrule
rule s1624(sum_count == 1624);
  total_sum <= total_sum + cache[1623];
endrule
rule s1625(sum_count == 1625);
  total_sum <= total_sum + cache[1624];
endrule
rule s1626(sum_count == 1626);
  total_sum <= total_sum + cache[1625];
endrule
rule s1627(sum_count == 1627);
  total_sum <= total_sum + cache[1626];
endrule
rule s1628(sum_count == 1628);
  total_sum <= total_sum + cache[1627];
endrule
rule s1629(sum_count == 1629);
  total_sum <= total_sum + cache[1628];
endrule
rule s1630(sum_count == 1630);
  total_sum <= total_sum + cache[1629];
endrule
rule s1631(sum_count == 1631);
  total_sum <= total_sum + cache[1630];
endrule
rule s1632(sum_count == 1632);
  total_sum <= total_sum + cache[1631];
endrule
rule s1633(sum_count == 1633);
  total_sum <= total_sum + cache[1632];
endrule
rule s1634(sum_count == 1634);
  total_sum <= total_sum + cache[1633];
endrule
rule s1635(sum_count == 1635);
  total_sum <= total_sum + cache[1634];
endrule
rule s1636(sum_count == 1636);
  total_sum <= total_sum + cache[1635];
endrule
rule s1637(sum_count == 1637);
  total_sum <= total_sum + cache[1636];
endrule
rule s1638(sum_count == 1638);
  total_sum <= total_sum + cache[1637];
endrule
rule s1639(sum_count == 1639);
  total_sum <= total_sum + cache[1638];
endrule
rule s1640(sum_count == 1640);
  total_sum <= total_sum + cache[1639];
endrule
rule s1641(sum_count == 1641);
  total_sum <= total_sum + cache[1640];
endrule
rule s1642(sum_count == 1642);
  total_sum <= total_sum + cache[1641];
endrule
rule s1643(sum_count == 1643);
  total_sum <= total_sum + cache[1642];
endrule
rule s1644(sum_count == 1644);
  total_sum <= total_sum + cache[1643];
endrule
rule s1645(sum_count == 1645);
  total_sum <= total_sum + cache[1644];
endrule
rule s1646(sum_count == 1646);
  total_sum <= total_sum + cache[1645];
endrule
rule s1647(sum_count == 1647);
  total_sum <= total_sum + cache[1646];
endrule
rule s1648(sum_count == 1648);
  total_sum <= total_sum + cache[1647];
endrule
rule s1649(sum_count == 1649);
  total_sum <= total_sum + cache[1648];
endrule
rule s1650(sum_count == 1650);
  total_sum <= total_sum + cache[1649];
endrule
rule s1651(sum_count == 1651);
  total_sum <= total_sum + cache[1650];
endrule
rule s1652(sum_count == 1652);
  total_sum <= total_sum + cache[1651];
endrule
rule s1653(sum_count == 1653);
  total_sum <= total_sum + cache[1652];
endrule
rule s1654(sum_count == 1654);
  total_sum <= total_sum + cache[1653];
endrule
rule s1655(sum_count == 1655);
  total_sum <= total_sum + cache[1654];
endrule
rule s1656(sum_count == 1656);
  total_sum <= total_sum + cache[1655];
endrule
rule s1657(sum_count == 1657);
  total_sum <= total_sum + cache[1656];
endrule
rule s1658(sum_count == 1658);
  total_sum <= total_sum + cache[1657];
endrule
rule s1659(sum_count == 1659);
  total_sum <= total_sum + cache[1658];
endrule
rule s1660(sum_count == 1660);
  total_sum <= total_sum + cache[1659];
endrule
rule s1661(sum_count == 1661);
  total_sum <= total_sum + cache[1660];
endrule
rule s1662(sum_count == 1662);
  total_sum <= total_sum + cache[1661];
endrule
rule s1663(sum_count == 1663);
  total_sum <= total_sum + cache[1662];
endrule
rule s1664(sum_count == 1664);
  total_sum <= total_sum + cache[1663];
endrule
rule s1665(sum_count == 1665);
  total_sum <= total_sum + cache[1664];
endrule
rule s1666(sum_count == 1666);
  total_sum <= total_sum + cache[1665];
endrule
rule s1667(sum_count == 1667);
  total_sum <= total_sum + cache[1666];
endrule
rule s1668(sum_count == 1668);
  total_sum <= total_sum + cache[1667];
endrule
rule s1669(sum_count == 1669);
  total_sum <= total_sum + cache[1668];
endrule
rule s1670(sum_count == 1670);
  total_sum <= total_sum + cache[1669];
endrule
rule s1671(sum_count == 1671);
  total_sum <= total_sum + cache[1670];
endrule
rule s1672(sum_count == 1672);
  total_sum <= total_sum + cache[1671];
endrule
rule s1673(sum_count == 1673);
  total_sum <= total_sum + cache[1672];
endrule
rule s1674(sum_count == 1674);
  total_sum <= total_sum + cache[1673];
endrule
rule s1675(sum_count == 1675);
  total_sum <= total_sum + cache[1674];
endrule
rule s1676(sum_count == 1676);
  total_sum <= total_sum + cache[1675];
endrule
rule s1677(sum_count == 1677);
  total_sum <= total_sum + cache[1676];
endrule
rule s1678(sum_count == 1678);
  total_sum <= total_sum + cache[1677];
endrule
rule s1679(sum_count == 1679);
  total_sum <= total_sum + cache[1678];
endrule
rule s1680(sum_count == 1680);
  total_sum <= total_sum + cache[1679];
endrule
rule s1681(sum_count == 1681);
  total_sum <= total_sum + cache[1680];
endrule
rule s1682(sum_count == 1682);
  total_sum <= total_sum + cache[1681];
endrule
rule s1683(sum_count == 1683);
  total_sum <= total_sum + cache[1682];
endrule
rule s1684(sum_count == 1684);
  total_sum <= total_sum + cache[1683];
endrule
rule s1685(sum_count == 1685);
  total_sum <= total_sum + cache[1684];
endrule
rule s1686(sum_count == 1686);
  total_sum <= total_sum + cache[1685];
endrule
rule s1687(sum_count == 1687);
  total_sum <= total_sum + cache[1686];
endrule
rule s1688(sum_count == 1688);
  total_sum <= total_sum + cache[1687];
endrule
rule s1689(sum_count == 1689);
  total_sum <= total_sum + cache[1688];
endrule
rule s1690(sum_count == 1690);
  total_sum <= total_sum + cache[1689];
endrule
rule s1691(sum_count == 1691);
  total_sum <= total_sum + cache[1690];
endrule
rule s1692(sum_count == 1692);
  total_sum <= total_sum + cache[1691];
endrule
rule s1693(sum_count == 1693);
  total_sum <= total_sum + cache[1692];
endrule
rule s1694(sum_count == 1694);
  total_sum <= total_sum + cache[1693];
endrule
rule s1695(sum_count == 1695);
  total_sum <= total_sum + cache[1694];
endrule
rule s1696(sum_count == 1696);
  total_sum <= total_sum + cache[1695];
endrule
rule s1697(sum_count == 1697);
  total_sum <= total_sum + cache[1696];
endrule
rule s1698(sum_count == 1698);
  total_sum <= total_sum + cache[1697];
endrule
rule s1699(sum_count == 1699);
  total_sum <= total_sum + cache[1698];
endrule
rule s1700(sum_count == 1700);
  total_sum <= total_sum + cache[1699];
endrule
rule s1701(sum_count == 1701);
  total_sum <= total_sum + cache[1700];
endrule
rule s1702(sum_count == 1702);
  total_sum <= total_sum + cache[1701];
endrule
rule s1703(sum_count == 1703);
  total_sum <= total_sum + cache[1702];
endrule
rule s1704(sum_count == 1704);
  total_sum <= total_sum + cache[1703];
endrule
rule s1705(sum_count == 1705);
  total_sum <= total_sum + cache[1704];
endrule
rule s1706(sum_count == 1706);
  total_sum <= total_sum + cache[1705];
endrule
rule s1707(sum_count == 1707);
  total_sum <= total_sum + cache[1706];
endrule
rule s1708(sum_count == 1708);
  total_sum <= total_sum + cache[1707];
endrule
rule s1709(sum_count == 1709);
  total_sum <= total_sum + cache[1708];
endrule
rule s1710(sum_count == 1710);
  total_sum <= total_sum + cache[1709];
endrule
rule s1711(sum_count == 1711);
  total_sum <= total_sum + cache[1710];
endrule
rule s1712(sum_count == 1712);
  total_sum <= total_sum + cache[1711];
endrule
rule s1713(sum_count == 1713);
  total_sum <= total_sum + cache[1712];
endrule
rule s1714(sum_count == 1714);
  total_sum <= total_sum + cache[1713];
endrule
rule s1715(sum_count == 1715);
  total_sum <= total_sum + cache[1714];
endrule
rule s1716(sum_count == 1716);
  total_sum <= total_sum + cache[1715];
endrule
rule s1717(sum_count == 1717);
  total_sum <= total_sum + cache[1716];
endrule
rule s1718(sum_count == 1718);
  total_sum <= total_sum + cache[1717];
endrule
rule s1719(sum_count == 1719);
  total_sum <= total_sum + cache[1718];
endrule
rule s1720(sum_count == 1720);
  total_sum <= total_sum + cache[1719];
endrule
rule s1721(sum_count == 1721);
  total_sum <= total_sum + cache[1720];
endrule
rule s1722(sum_count == 1722);
  total_sum <= total_sum + cache[1721];
endrule
rule s1723(sum_count == 1723);
  total_sum <= total_sum + cache[1722];
endrule
rule s1724(sum_count == 1724);
  total_sum <= total_sum + cache[1723];
endrule
rule s1725(sum_count == 1725);
  total_sum <= total_sum + cache[1724];
endrule
rule s1726(sum_count == 1726);
  total_sum <= total_sum + cache[1725];
endrule
rule s1727(sum_count == 1727);
  total_sum <= total_sum + cache[1726];
endrule
rule s1728(sum_count == 1728);
  total_sum <= total_sum + cache[1727];
endrule
rule s1729(sum_count == 1729);
  total_sum <= total_sum + cache[1728];
endrule
rule s1730(sum_count == 1730);
  total_sum <= total_sum + cache[1729];
endrule
rule s1731(sum_count == 1731);
  total_sum <= total_sum + cache[1730];
endrule
rule s1732(sum_count == 1732);
  total_sum <= total_sum + cache[1731];
endrule
rule s1733(sum_count == 1733);
  total_sum <= total_sum + cache[1732];
endrule
rule s1734(sum_count == 1734);
  total_sum <= total_sum + cache[1733];
endrule
rule s1735(sum_count == 1735);
  total_sum <= total_sum + cache[1734];
endrule
rule s1736(sum_count == 1736);
  total_sum <= total_sum + cache[1735];
endrule
rule s1737(sum_count == 1737);
  total_sum <= total_sum + cache[1736];
endrule
rule s1738(sum_count == 1738);
  total_sum <= total_sum + cache[1737];
endrule
rule s1739(sum_count == 1739);
  total_sum <= total_sum + cache[1738];
endrule
rule s1740(sum_count == 1740);
  total_sum <= total_sum + cache[1739];
endrule
rule s1741(sum_count == 1741);
  total_sum <= total_sum + cache[1740];
endrule
rule s1742(sum_count == 1742);
  total_sum <= total_sum + cache[1741];
endrule
rule s1743(sum_count == 1743);
  total_sum <= total_sum + cache[1742];
endrule
rule s1744(sum_count == 1744);
  total_sum <= total_sum + cache[1743];
endrule
rule s1745(sum_count == 1745);
  total_sum <= total_sum + cache[1744];
endrule
rule s1746(sum_count == 1746);
  total_sum <= total_sum + cache[1745];
endrule
rule s1747(sum_count == 1747);
  total_sum <= total_sum + cache[1746];
endrule
rule s1748(sum_count == 1748);
  total_sum <= total_sum + cache[1747];
endrule
rule s1749(sum_count == 1749);
  total_sum <= total_sum + cache[1748];
endrule
rule s1750(sum_count == 1750);
  total_sum <= total_sum + cache[1749];
endrule
rule s1751(sum_count == 1751);
  total_sum <= total_sum + cache[1750];
endrule
rule s1752(sum_count == 1752);
  total_sum <= total_sum + cache[1751];
endrule
rule s1753(sum_count == 1753);
  total_sum <= total_sum + cache[1752];
endrule
rule s1754(sum_count == 1754);
  total_sum <= total_sum + cache[1753];
endrule
rule s1755(sum_count == 1755);
  total_sum <= total_sum + cache[1754];
endrule
rule s1756(sum_count == 1756);
  total_sum <= total_sum + cache[1755];
endrule
rule s1757(sum_count == 1757);
  total_sum <= total_sum + cache[1756];
endrule
rule s1758(sum_count == 1758);
  total_sum <= total_sum + cache[1757];
endrule
rule s1759(sum_count == 1759);
  total_sum <= total_sum + cache[1758];
endrule
rule s1760(sum_count == 1760);
  total_sum <= total_sum + cache[1759];
endrule
rule s1761(sum_count == 1761);
  total_sum <= total_sum + cache[1760];
endrule
rule s1762(sum_count == 1762);
  total_sum <= total_sum + cache[1761];
endrule
rule s1763(sum_count == 1763);
  total_sum <= total_sum + cache[1762];
endrule
rule s1764(sum_count == 1764);
  total_sum <= total_sum + cache[1763];
endrule
rule s1765(sum_count == 1765);
  total_sum <= total_sum + cache[1764];
endrule
rule s1766(sum_count == 1766);
  total_sum <= total_sum + cache[1765];
endrule
rule s1767(sum_count == 1767);
  total_sum <= total_sum + cache[1766];
endrule
rule s1768(sum_count == 1768);
  total_sum <= total_sum + cache[1767];
endrule
rule s1769(sum_count == 1769);
  total_sum <= total_sum + cache[1768];
endrule
rule s1770(sum_count == 1770);
  total_sum <= total_sum + cache[1769];
endrule
rule s1771(sum_count == 1771);
  total_sum <= total_sum + cache[1770];
endrule
rule s1772(sum_count == 1772);
  total_sum <= total_sum + cache[1771];
endrule
rule s1773(sum_count == 1773);
  total_sum <= total_sum + cache[1772];
endrule
rule s1774(sum_count == 1774);
  total_sum <= total_sum + cache[1773];
endrule
rule s1775(sum_count == 1775);
  total_sum <= total_sum + cache[1774];
endrule
rule s1776(sum_count == 1776);
  total_sum <= total_sum + cache[1775];
endrule
rule s1777(sum_count == 1777);
  total_sum <= total_sum + cache[1776];
endrule
rule s1778(sum_count == 1778);
  total_sum <= total_sum + cache[1777];
endrule
rule s1779(sum_count == 1779);
  total_sum <= total_sum + cache[1778];
endrule
rule s1780(sum_count == 1780);
  total_sum <= total_sum + cache[1779];
endrule
rule s1781(sum_count == 1781);
  total_sum <= total_sum + cache[1780];
endrule
rule s1782(sum_count == 1782);
  total_sum <= total_sum + cache[1781];
endrule
rule s1783(sum_count == 1783);
  total_sum <= total_sum + cache[1782];
endrule
rule s1784(sum_count == 1784);
  total_sum <= total_sum + cache[1783];
endrule
rule s1785(sum_count == 1785);
  total_sum <= total_sum + cache[1784];
endrule
rule s1786(sum_count == 1786);
  total_sum <= total_sum + cache[1785];
endrule
rule s1787(sum_count == 1787);
  total_sum <= total_sum + cache[1786];
endrule
rule s1788(sum_count == 1788);
  total_sum <= total_sum + cache[1787];
endrule
rule s1789(sum_count == 1789);
  total_sum <= total_sum + cache[1788];
endrule
rule s1790(sum_count == 1790);
  total_sum <= total_sum + cache[1789];
endrule
rule s1791(sum_count == 1791);
  total_sum <= total_sum + cache[1790];
endrule
rule s1792(sum_count == 1792);
  total_sum <= total_sum + cache[1791];
endrule
rule s1793(sum_count == 1793);
  total_sum <= total_sum + cache[1792];
endrule
rule s1794(sum_count == 1794);
  total_sum <= total_sum + cache[1793];
endrule
rule s1795(sum_count == 1795);
  total_sum <= total_sum + cache[1794];
endrule
rule s1796(sum_count == 1796);
  total_sum <= total_sum + cache[1795];
endrule
rule s1797(sum_count == 1797);
  total_sum <= total_sum + cache[1796];
endrule
rule s1798(sum_count == 1798);
  total_sum <= total_sum + cache[1797];
endrule
rule s1799(sum_count == 1799);
  total_sum <= total_sum + cache[1798];
endrule
rule s1800(sum_count == 1800);
  total_sum <= total_sum + cache[1799];
endrule
rule s1801(sum_count == 1801);
  total_sum <= total_sum + cache[1800];
endrule
rule s1802(sum_count == 1802);
  total_sum <= total_sum + cache[1801];
endrule
rule s1803(sum_count == 1803);
  total_sum <= total_sum + cache[1802];
endrule
rule s1804(sum_count == 1804);
  total_sum <= total_sum + cache[1803];
endrule
rule s1805(sum_count == 1805);
  total_sum <= total_sum + cache[1804];
endrule
rule s1806(sum_count == 1806);
  total_sum <= total_sum + cache[1805];
endrule
rule s1807(sum_count == 1807);
  total_sum <= total_sum + cache[1806];
endrule
rule s1808(sum_count == 1808);
  total_sum <= total_sum + cache[1807];
endrule
rule s1809(sum_count == 1809);
  total_sum <= total_sum + cache[1808];
endrule
rule s1810(sum_count == 1810);
  total_sum <= total_sum + cache[1809];
endrule
rule s1811(sum_count == 1811);
  total_sum <= total_sum + cache[1810];
endrule
rule s1812(sum_count == 1812);
  total_sum <= total_sum + cache[1811];
endrule
rule s1813(sum_count == 1813);
  total_sum <= total_sum + cache[1812];
endrule
rule s1814(sum_count == 1814);
  total_sum <= total_sum + cache[1813];
endrule
rule s1815(sum_count == 1815);
  total_sum <= total_sum + cache[1814];
endrule
rule s1816(sum_count == 1816);
  total_sum <= total_sum + cache[1815];
endrule
rule s1817(sum_count == 1817);
  total_sum <= total_sum + cache[1816];
endrule
rule s1818(sum_count == 1818);
  total_sum <= total_sum + cache[1817];
endrule
rule s1819(sum_count == 1819);
  total_sum <= total_sum + cache[1818];
endrule
rule s1820(sum_count == 1820);
  total_sum <= total_sum + cache[1819];
endrule
rule s1821(sum_count == 1821);
  total_sum <= total_sum + cache[1820];
endrule
rule s1822(sum_count == 1822);
  total_sum <= total_sum + cache[1821];
endrule
rule s1823(sum_count == 1823);
  total_sum <= total_sum + cache[1822];
endrule
rule s1824(sum_count == 1824);
  total_sum <= total_sum + cache[1823];
endrule
rule s1825(sum_count == 1825);
  total_sum <= total_sum + cache[1824];
endrule
rule s1826(sum_count == 1826);
  total_sum <= total_sum + cache[1825];
endrule
rule s1827(sum_count == 1827);
  total_sum <= total_sum + cache[1826];
endrule
rule s1828(sum_count == 1828);
  total_sum <= total_sum + cache[1827];
endrule
rule s1829(sum_count == 1829);
  total_sum <= total_sum + cache[1828];
endrule
rule s1830(sum_count == 1830);
  total_sum <= total_sum + cache[1829];
endrule
rule s1831(sum_count == 1831);
  total_sum <= total_sum + cache[1830];
endrule
rule s1832(sum_count == 1832);
  total_sum <= total_sum + cache[1831];
endrule
rule s1833(sum_count == 1833);
  total_sum <= total_sum + cache[1832];
endrule
rule s1834(sum_count == 1834);
  total_sum <= total_sum + cache[1833];
endrule
rule s1835(sum_count == 1835);
  total_sum <= total_sum + cache[1834];
endrule
rule s1836(sum_count == 1836);
  total_sum <= total_sum + cache[1835];
endrule
rule s1837(sum_count == 1837);
  total_sum <= total_sum + cache[1836];
endrule
rule s1838(sum_count == 1838);
  total_sum <= total_sum + cache[1837];
endrule
rule s1839(sum_count == 1839);
  total_sum <= total_sum + cache[1838];
endrule
rule s1840(sum_count == 1840);
  total_sum <= total_sum + cache[1839];
endrule
rule s1841(sum_count == 1841);
  total_sum <= total_sum + cache[1840];
endrule
rule s1842(sum_count == 1842);
  total_sum <= total_sum + cache[1841];
endrule
rule s1843(sum_count == 1843);
  total_sum <= total_sum + cache[1842];
endrule
rule s1844(sum_count == 1844);
  total_sum <= total_sum + cache[1843];
endrule
rule s1845(sum_count == 1845);
  total_sum <= total_sum + cache[1844];
endrule
rule s1846(sum_count == 1846);
  total_sum <= total_sum + cache[1845];
endrule
rule s1847(sum_count == 1847);
  total_sum <= total_sum + cache[1846];
endrule
rule s1848(sum_count == 1848);
  total_sum <= total_sum + cache[1847];
endrule
rule s1849(sum_count == 1849);
  total_sum <= total_sum + cache[1848];
endrule
rule s1850(sum_count == 1850);
  total_sum <= total_sum + cache[1849];
endrule
rule s1851(sum_count == 1851);
  total_sum <= total_sum + cache[1850];
endrule
rule s1852(sum_count == 1852);
  total_sum <= total_sum + cache[1851];
endrule
rule s1853(sum_count == 1853);
  total_sum <= total_sum + cache[1852];
endrule
rule s1854(sum_count == 1854);
  total_sum <= total_sum + cache[1853];
endrule
rule s1855(sum_count == 1855);
  total_sum <= total_sum + cache[1854];
endrule
rule s1856(sum_count == 1856);
  total_sum <= total_sum + cache[1855];
endrule
rule s1857(sum_count == 1857);
  total_sum <= total_sum + cache[1856];
endrule
rule s1858(sum_count == 1858);
  total_sum <= total_sum + cache[1857];
endrule
rule s1859(sum_count == 1859);
  total_sum <= total_sum + cache[1858];
endrule
rule s1860(sum_count == 1860);
  total_sum <= total_sum + cache[1859];
endrule
rule s1861(sum_count == 1861);
  total_sum <= total_sum + cache[1860];
endrule
rule s1862(sum_count == 1862);
  total_sum <= total_sum + cache[1861];
endrule
rule s1863(sum_count == 1863);
  total_sum <= total_sum + cache[1862];
endrule
rule s1864(sum_count == 1864);
  total_sum <= total_sum + cache[1863];
endrule
rule s1865(sum_count == 1865);
  total_sum <= total_sum + cache[1864];
endrule
rule s1866(sum_count == 1866);
  total_sum <= total_sum + cache[1865];
endrule
rule s1867(sum_count == 1867);
  total_sum <= total_sum + cache[1866];
endrule
rule s1868(sum_count == 1868);
  total_sum <= total_sum + cache[1867];
endrule
rule s1869(sum_count == 1869);
  total_sum <= total_sum + cache[1868];
endrule
rule s1870(sum_count == 1870);
  total_sum <= total_sum + cache[1869];
endrule
rule s1871(sum_count == 1871);
  total_sum <= total_sum + cache[1870];
endrule
rule s1872(sum_count == 1872);
  total_sum <= total_sum + cache[1871];
endrule
rule s1873(sum_count == 1873);
  total_sum <= total_sum + cache[1872];
endrule
rule s1874(sum_count == 1874);
  total_sum <= total_sum + cache[1873];
endrule
rule s1875(sum_count == 1875);
  total_sum <= total_sum + cache[1874];
endrule
rule s1876(sum_count == 1876);
  total_sum <= total_sum + cache[1875];
endrule
rule s1877(sum_count == 1877);
  total_sum <= total_sum + cache[1876];
endrule
rule s1878(sum_count == 1878);
  total_sum <= total_sum + cache[1877];
endrule
rule s1879(sum_count == 1879);
  total_sum <= total_sum + cache[1878];
endrule
rule s1880(sum_count == 1880);
  total_sum <= total_sum + cache[1879];
endrule
rule s1881(sum_count == 1881);
  total_sum <= total_sum + cache[1880];
endrule
rule s1882(sum_count == 1882);
  total_sum <= total_sum + cache[1881];
endrule
rule s1883(sum_count == 1883);
  total_sum <= total_sum + cache[1882];
endrule
rule s1884(sum_count == 1884);
  total_sum <= total_sum + cache[1883];
endrule
rule s1885(sum_count == 1885);
  total_sum <= total_sum + cache[1884];
endrule
rule s1886(sum_count == 1886);
  total_sum <= total_sum + cache[1885];
endrule
rule s1887(sum_count == 1887);
  total_sum <= total_sum + cache[1886];
endrule
rule s1888(sum_count == 1888);
  total_sum <= total_sum + cache[1887];
endrule
rule s1889(sum_count == 1889);
  total_sum <= total_sum + cache[1888];
endrule
rule s1890(sum_count == 1890);
  total_sum <= total_sum + cache[1889];
endrule
rule s1891(sum_count == 1891);
  total_sum <= total_sum + cache[1890];
endrule
rule s1892(sum_count == 1892);
  total_sum <= total_sum + cache[1891];
endrule
rule s1893(sum_count == 1893);
  total_sum <= total_sum + cache[1892];
endrule
rule s1894(sum_count == 1894);
  total_sum <= total_sum + cache[1893];
endrule
rule s1895(sum_count == 1895);
  total_sum <= total_sum + cache[1894];
endrule
rule s1896(sum_count == 1896);
  total_sum <= total_sum + cache[1895];
endrule
rule s1897(sum_count == 1897);
  total_sum <= total_sum + cache[1896];
endrule
rule s1898(sum_count == 1898);
  total_sum <= total_sum + cache[1897];
endrule
rule s1899(sum_count == 1899);
  total_sum <= total_sum + cache[1898];
endrule
rule s1900(sum_count == 1900);
  total_sum <= total_sum + cache[1899];
endrule
rule s1901(sum_count == 1901);
  total_sum <= total_sum + cache[1900];
endrule
rule s1902(sum_count == 1902);
  total_sum <= total_sum + cache[1901];
endrule
rule s1903(sum_count == 1903);
  total_sum <= total_sum + cache[1902];
endrule
rule s1904(sum_count == 1904);
  total_sum <= total_sum + cache[1903];
endrule
rule s1905(sum_count == 1905);
  total_sum <= total_sum + cache[1904];
endrule
rule s1906(sum_count == 1906);
  total_sum <= total_sum + cache[1905];
endrule
rule s1907(sum_count == 1907);
  total_sum <= total_sum + cache[1906];
endrule
rule s1908(sum_count == 1908);
  total_sum <= total_sum + cache[1907];
endrule
rule s1909(sum_count == 1909);
  total_sum <= total_sum + cache[1908];
endrule
rule s1910(sum_count == 1910);
  total_sum <= total_sum + cache[1909];
endrule
rule s1911(sum_count == 1911);
  total_sum <= total_sum + cache[1910];
endrule
rule s1912(sum_count == 1912);
  total_sum <= total_sum + cache[1911];
endrule
rule s1913(sum_count == 1913);
  total_sum <= total_sum + cache[1912];
endrule
rule s1914(sum_count == 1914);
  total_sum <= total_sum + cache[1913];
endrule
rule s1915(sum_count == 1915);
  total_sum <= total_sum + cache[1914];
endrule
rule s1916(sum_count == 1916);
  total_sum <= total_sum + cache[1915];
endrule
rule s1917(sum_count == 1917);
  total_sum <= total_sum + cache[1916];
endrule
rule s1918(sum_count == 1918);
  total_sum <= total_sum + cache[1917];
endrule
rule s1919(sum_count == 1919);
  total_sum <= total_sum + cache[1918];
endrule
rule s1920(sum_count == 1920);
  total_sum <= total_sum + cache[1919];
endrule
rule s1921(sum_count == 1921);
  total_sum <= total_sum + cache[1920];
endrule
rule s1922(sum_count == 1922);
  total_sum <= total_sum + cache[1921];
endrule
rule s1923(sum_count == 1923);
  total_sum <= total_sum + cache[1922];
endrule
rule s1924(sum_count == 1924);
  total_sum <= total_sum + cache[1923];
endrule
rule s1925(sum_count == 1925);
  total_sum <= total_sum + cache[1924];
endrule
rule s1926(sum_count == 1926);
  total_sum <= total_sum + cache[1925];
endrule
rule s1927(sum_count == 1927);
  total_sum <= total_sum + cache[1926];
endrule
rule s1928(sum_count == 1928);
  total_sum <= total_sum + cache[1927];
endrule
rule s1929(sum_count == 1929);
  total_sum <= total_sum + cache[1928];
endrule
rule s1930(sum_count == 1930);
  total_sum <= total_sum + cache[1929];
endrule
rule s1931(sum_count == 1931);
  total_sum <= total_sum + cache[1930];
endrule
rule s1932(sum_count == 1932);
  total_sum <= total_sum + cache[1931];
endrule
rule s1933(sum_count == 1933);
  total_sum <= total_sum + cache[1932];
endrule
rule s1934(sum_count == 1934);
  total_sum <= total_sum + cache[1933];
endrule
rule s1935(sum_count == 1935);
  total_sum <= total_sum + cache[1934];
endrule
rule s1936(sum_count == 1936);
  total_sum <= total_sum + cache[1935];
endrule
rule s1937(sum_count == 1937);
  total_sum <= total_sum + cache[1936];
endrule
rule s1938(sum_count == 1938);
  total_sum <= total_sum + cache[1937];
endrule
rule s1939(sum_count == 1939);
  total_sum <= total_sum + cache[1938];
endrule
rule s1940(sum_count == 1940);
  total_sum <= total_sum + cache[1939];
endrule
rule s1941(sum_count == 1941);
  total_sum <= total_sum + cache[1940];
endrule
rule s1942(sum_count == 1942);
  total_sum <= total_sum + cache[1941];
endrule
rule s1943(sum_count == 1943);
  total_sum <= total_sum + cache[1942];
endrule
rule s1944(sum_count == 1944);
  total_sum <= total_sum + cache[1943];
endrule
rule s1945(sum_count == 1945);
  total_sum <= total_sum + cache[1944];
endrule
rule s1946(sum_count == 1946);
  total_sum <= total_sum + cache[1945];
endrule
rule s1947(sum_count == 1947);
  total_sum <= total_sum + cache[1946];
endrule
rule s1948(sum_count == 1948);
  total_sum <= total_sum + cache[1947];
endrule
rule s1949(sum_count == 1949);
  total_sum <= total_sum + cache[1948];
endrule
rule s1950(sum_count == 1950);
  total_sum <= total_sum + cache[1949];
endrule
rule s1951(sum_count == 1951);
  total_sum <= total_sum + cache[1950];
endrule
rule s1952(sum_count == 1952);
  total_sum <= total_sum + cache[1951];
endrule
rule s1953(sum_count == 1953);
  total_sum <= total_sum + cache[1952];
endrule
rule s1954(sum_count == 1954);
  total_sum <= total_sum + cache[1953];
endrule
rule s1955(sum_count == 1955);
  total_sum <= total_sum + cache[1954];
endrule
rule s1956(sum_count == 1956);
  total_sum <= total_sum + cache[1955];
endrule
rule s1957(sum_count == 1957);
  total_sum <= total_sum + cache[1956];
endrule
rule s1958(sum_count == 1958);
  total_sum <= total_sum + cache[1957];
endrule
rule s1959(sum_count == 1959);
  total_sum <= total_sum + cache[1958];
endrule
rule s1960(sum_count == 1960);
  total_sum <= total_sum + cache[1959];
endrule
rule s1961(sum_count == 1961);
  total_sum <= total_sum + cache[1960];
endrule
rule s1962(sum_count == 1962);
  total_sum <= total_sum + cache[1961];
endrule
rule s1963(sum_count == 1963);
  total_sum <= total_sum + cache[1962];
endrule
rule s1964(sum_count == 1964);
  total_sum <= total_sum + cache[1963];
endrule
rule s1965(sum_count == 1965);
  total_sum <= total_sum + cache[1964];
endrule
rule s1966(sum_count == 1966);
  total_sum <= total_sum + cache[1965];
endrule
rule s1967(sum_count == 1967);
  total_sum <= total_sum + cache[1966];
endrule
rule s1968(sum_count == 1968);
  total_sum <= total_sum + cache[1967];
endrule
rule s1969(sum_count == 1969);
  total_sum <= total_sum + cache[1968];
endrule
rule s1970(sum_count == 1970);
  total_sum <= total_sum + cache[1969];
endrule
rule s1971(sum_count == 1971);
  total_sum <= total_sum + cache[1970];
endrule
rule s1972(sum_count == 1972);
  total_sum <= total_sum + cache[1971];
endrule
rule s1973(sum_count == 1973);
  total_sum <= total_sum + cache[1972];
endrule
rule s1974(sum_count == 1974);
  total_sum <= total_sum + cache[1973];
endrule
rule s1975(sum_count == 1975);
  total_sum <= total_sum + cache[1974];
endrule
rule s1976(sum_count == 1976);
  total_sum <= total_sum + cache[1975];
endrule
rule s1977(sum_count == 1977);
  total_sum <= total_sum + cache[1976];
endrule
rule s1978(sum_count == 1978);
  total_sum <= total_sum + cache[1977];
endrule
rule s1979(sum_count == 1979);
  total_sum <= total_sum + cache[1978];
endrule
rule s1980(sum_count == 1980);
  total_sum <= total_sum + cache[1979];
endrule
rule s1981(sum_count == 1981);
  total_sum <= total_sum + cache[1980];
endrule
rule s1982(sum_count == 1982);
  total_sum <= total_sum + cache[1981];
endrule
rule s1983(sum_count == 1983);
  total_sum <= total_sum + cache[1982];
endrule
rule s1984(sum_count == 1984);
  total_sum <= total_sum + cache[1983];
endrule
rule s1985(sum_count == 1985);
  total_sum <= total_sum + cache[1984];
endrule
rule s1986(sum_count == 1986);
  total_sum <= total_sum + cache[1985];
endrule
rule s1987(sum_count == 1987);
  total_sum <= total_sum + cache[1986];
endrule
rule s1988(sum_count == 1988);
  total_sum <= total_sum + cache[1987];
endrule
rule s1989(sum_count == 1989);
  total_sum <= total_sum + cache[1988];
endrule
rule s1990(sum_count == 1990);
  total_sum <= total_sum + cache[1989];
endrule
rule s1991(sum_count == 1991);
  total_sum <= total_sum + cache[1990];
endrule
rule s1992(sum_count == 1992);
  total_sum <= total_sum + cache[1991];
endrule
rule s1993(sum_count == 1993);
  total_sum <= total_sum + cache[1992];
endrule
rule s1994(sum_count == 1994);
  total_sum <= total_sum + cache[1993];
endrule
rule s1995(sum_count == 1995);
  total_sum <= total_sum + cache[1994];
endrule
rule s1996(sum_count == 1996);
  total_sum <= total_sum + cache[1995];
endrule
rule s1997(sum_count == 1997);
  total_sum <= total_sum + cache[1996];
endrule
rule s1998(sum_count == 1998);
  total_sum <= total_sum + cache[1997];
endrule
rule s1999(sum_count == 1999);
  total_sum <= total_sum + cache[1998];
endrule
rule s2000(sum_count == 2000);
  total_sum <= total_sum + cache[1999];
endrule
rule s2001(sum_count == 2001);
  total_sum <= total_sum + cache[2000];
endrule
rule s2002(sum_count == 2002);
  total_sum <= total_sum + cache[2001];
endrule
rule s2003(sum_count == 2003);
  total_sum <= total_sum + cache[2002];
endrule
rule s2004(sum_count == 2004);
  total_sum <= total_sum + cache[2003];
endrule
rule s2005(sum_count == 2005);
  total_sum <= total_sum + cache[2004];
endrule
rule s2006(sum_count == 2006);
  total_sum <= total_sum + cache[2005];
endrule
rule s2007(sum_count == 2007);
  total_sum <= total_sum + cache[2006];
endrule
rule s2008(sum_count == 2008);
  total_sum <= total_sum + cache[2007];
endrule
rule s2009(sum_count == 2009);
  total_sum <= total_sum + cache[2008];
endrule
rule s2010(sum_count == 2010);
  total_sum <= total_sum + cache[2009];
endrule
rule s2011(sum_count == 2011);
  total_sum <= total_sum + cache[2010];
endrule
rule s2012(sum_count == 2012);
  total_sum <= total_sum + cache[2011];
endrule
rule s2013(sum_count == 2013);
  total_sum <= total_sum + cache[2012];
endrule
rule s2014(sum_count == 2014);
  total_sum <= total_sum + cache[2013];
endrule
rule s2015(sum_count == 2015);
  total_sum <= total_sum + cache[2014];
endrule
rule s2016(sum_count == 2016);
  total_sum <= total_sum + cache[2015];
endrule
rule s2017(sum_count == 2017);
  total_sum <= total_sum + cache[2016];
endrule
rule s2018(sum_count == 2018);
  total_sum <= total_sum + cache[2017];
endrule
rule s2019(sum_count == 2019);
  total_sum <= total_sum + cache[2018];
endrule
rule s2020(sum_count == 2020);
  total_sum <= total_sum + cache[2019];
endrule
rule s2021(sum_count == 2021);
  total_sum <= total_sum + cache[2020];
endrule
rule s2022(sum_count == 2022);
  total_sum <= total_sum + cache[2021];
endrule
rule s2023(sum_count == 2023);
  total_sum <= total_sum + cache[2022];
endrule
rule s2024(sum_count == 2024);
  total_sum <= total_sum + cache[2023];
endrule
rule s2025(sum_count == 2025);
  total_sum <= total_sum + cache[2024];
endrule
rule s2026(sum_count == 2026);
  total_sum <= total_sum + cache[2025];
endrule
rule s2027(sum_count == 2027);
  total_sum <= total_sum + cache[2026];
endrule
rule s2028(sum_count == 2028);
  total_sum <= total_sum + cache[2027];
endrule
rule s2029(sum_count == 2029);
  total_sum <= total_sum + cache[2028];
endrule
rule s2030(sum_count == 2030);
  total_sum <= total_sum + cache[2029];
endrule
rule s2031(sum_count == 2031);
  total_sum <= total_sum + cache[2030];
endrule
rule s2032(sum_count == 2032);
  total_sum <= total_sum + cache[2031];
endrule
rule s2033(sum_count == 2033);
  total_sum <= total_sum + cache[2032];
endrule
rule s2034(sum_count == 2034);
  total_sum <= total_sum + cache[2033];
endrule
rule s2035(sum_count == 2035);
  total_sum <= total_sum + cache[2034];
endrule
rule s2036(sum_count == 2036);
  total_sum <= total_sum + cache[2035];
endrule
rule s2037(sum_count == 2037);
  total_sum <= total_sum + cache[2036];
endrule
rule s2038(sum_count == 2038);
  total_sum <= total_sum + cache[2037];
endrule
rule s2039(sum_count == 2039);
  total_sum <= total_sum + cache[2038];
endrule
rule s2040(sum_count == 2040);
  total_sum <= total_sum + cache[2039];
endrule
rule s2041(sum_count == 2041);
  total_sum <= total_sum + cache[2040];
endrule
rule s2042(sum_count == 2042);
  total_sum <= total_sum + cache[2041];
endrule
rule s2043(sum_count == 2043);
  total_sum <= total_sum + cache[2042];
endrule
rule s2044(sum_count == 2044);
  total_sum <= total_sum + cache[2043];
endrule
rule s2045(sum_count == 2045);
  total_sum <= total_sum + cache[2044];
endrule
rule s2046(sum_count == 2046);
  total_sum <= total_sum + cache[2045];
endrule
rule s2047(sum_count == 2047);
  total_sum <= total_sum + cache[2046];
endrule
rule s2048(sum_count == 2048);
  total_sum <= total_sum + cache[2047];
endrule
rule s2049(sum_count == 2049);
  total_sum <= total_sum + cache[2048];
endrule
rule s2050(sum_count == 2050);
  total_sum <= total_sum + cache[2049];
endrule
rule s2051(sum_count == 2051);
  total_sum <= total_sum + cache[2050];
endrule
rule s2052(sum_count == 2052);
  total_sum <= total_sum + cache[2051];
endrule
rule s2053(sum_count == 2053);
  total_sum <= total_sum + cache[2052];
endrule
rule s2054(sum_count == 2054);
  total_sum <= total_sum + cache[2053];
endrule
rule s2055(sum_count == 2055);
  total_sum <= total_sum + cache[2054];
endrule
rule s2056(sum_count == 2056);
  total_sum <= total_sum + cache[2055];
endrule
rule s2057(sum_count == 2057);
  total_sum <= total_sum + cache[2056];
endrule
rule s2058(sum_count == 2058);
  total_sum <= total_sum + cache[2057];
endrule
rule s2059(sum_count == 2059);
  total_sum <= total_sum + cache[2058];
endrule
rule s2060(sum_count == 2060);
  total_sum <= total_sum + cache[2059];
endrule
rule s2061(sum_count == 2061);
  total_sum <= total_sum + cache[2060];
endrule
rule s2062(sum_count == 2062);
  total_sum <= total_sum + cache[2061];
endrule
rule s2063(sum_count == 2063);
  total_sum <= total_sum + cache[2062];
endrule
rule s2064(sum_count == 2064);
  total_sum <= total_sum + cache[2063];
endrule
rule s2065(sum_count == 2065);
  total_sum <= total_sum + cache[2064];
endrule
rule s2066(sum_count == 2066);
  total_sum <= total_sum + cache[2065];
endrule
rule s2067(sum_count == 2067);
  total_sum <= total_sum + cache[2066];
endrule
rule s2068(sum_count == 2068);
  total_sum <= total_sum + cache[2067];
endrule
rule s2069(sum_count == 2069);
  total_sum <= total_sum + cache[2068];
endrule
rule s2070(sum_count == 2070);
  total_sum <= total_sum + cache[2069];
endrule
rule s2071(sum_count == 2071);
  total_sum <= total_sum + cache[2070];
endrule
rule s2072(sum_count == 2072);
  total_sum <= total_sum + cache[2071];
endrule
rule s2073(sum_count == 2073);
  total_sum <= total_sum + cache[2072];
endrule
rule s2074(sum_count == 2074);
  total_sum <= total_sum + cache[2073];
endrule
rule s2075(sum_count == 2075);
  total_sum <= total_sum + cache[2074];
endrule
rule s2076(sum_count == 2076);
  total_sum <= total_sum + cache[2075];
endrule
rule s2077(sum_count == 2077);
  total_sum <= total_sum + cache[2076];
endrule
rule s2078(sum_count == 2078);
  total_sum <= total_sum + cache[2077];
endrule
rule s2079(sum_count == 2079);
  total_sum <= total_sum + cache[2078];
endrule
rule s2080(sum_count == 2080);
  total_sum <= total_sum + cache[2079];
endrule
rule s2081(sum_count == 2081);
  total_sum <= total_sum + cache[2080];
endrule
rule s2082(sum_count == 2082);
  total_sum <= total_sum + cache[2081];
endrule
rule s2083(sum_count == 2083);
  total_sum <= total_sum + cache[2082];
endrule
rule s2084(sum_count == 2084);
  total_sum <= total_sum + cache[2083];
endrule
rule s2085(sum_count == 2085);
  total_sum <= total_sum + cache[2084];
endrule
rule s2086(sum_count == 2086);
  total_sum <= total_sum + cache[2085];
endrule
rule s2087(sum_count == 2087);
  total_sum <= total_sum + cache[2086];
endrule
rule s2088(sum_count == 2088);
  total_sum <= total_sum + cache[2087];
endrule
rule s2089(sum_count == 2089);
  total_sum <= total_sum + cache[2088];
endrule
rule s2090(sum_count == 2090);
  total_sum <= total_sum + cache[2089];
endrule
rule s2091(sum_count == 2091);
  total_sum <= total_sum + cache[2090];
endrule
rule s2092(sum_count == 2092);
  total_sum <= total_sum + cache[2091];
endrule
rule s2093(sum_count == 2093);
  total_sum <= total_sum + cache[2092];
endrule
rule s2094(sum_count == 2094);
  total_sum <= total_sum + cache[2093];
endrule
rule s2095(sum_count == 2095);
  total_sum <= total_sum + cache[2094];
endrule
rule s2096(sum_count == 2096);
  total_sum <= total_sum + cache[2095];
endrule
rule s2097(sum_count == 2097);
  total_sum <= total_sum + cache[2096];
endrule
rule s2098(sum_count == 2098);
  total_sum <= total_sum + cache[2097];
endrule
rule s2099(sum_count == 2099);
  total_sum <= total_sum + cache[2098];
endrule
rule s2100(sum_count == 2100);
  total_sum <= total_sum + cache[2099];
endrule
rule s2101(sum_count == 2101);
  total_sum <= total_sum + cache[2100];
endrule
rule s2102(sum_count == 2102);
  total_sum <= total_sum + cache[2101];
endrule
rule s2103(sum_count == 2103);
  total_sum <= total_sum + cache[2102];
endrule
rule s2104(sum_count == 2104);
  total_sum <= total_sum + cache[2103];
endrule
rule s2105(sum_count == 2105);
  total_sum <= total_sum + cache[2104];
endrule
rule s2106(sum_count == 2106);
  total_sum <= total_sum + cache[2105];
endrule
rule s2107(sum_count == 2107);
  total_sum <= total_sum + cache[2106];
endrule
rule s2108(sum_count == 2108);
  total_sum <= total_sum + cache[2107];
endrule
rule s2109(sum_count == 2109);
  total_sum <= total_sum + cache[2108];
endrule
rule s2110(sum_count == 2110);
  total_sum <= total_sum + cache[2109];
endrule
rule s2111(sum_count == 2111);
  total_sum <= total_sum + cache[2110];
endrule
rule s2112(sum_count == 2112);
  total_sum <= total_sum + cache[2111];
endrule
rule s2113(sum_count == 2113);
  total_sum <= total_sum + cache[2112];
endrule
rule s2114(sum_count == 2114);
  total_sum <= total_sum + cache[2113];
endrule
rule s2115(sum_count == 2115);
  total_sum <= total_sum + cache[2114];
endrule
rule s2116(sum_count == 2116);
  total_sum <= total_sum + cache[2115];
endrule
rule s2117(sum_count == 2117);
  total_sum <= total_sum + cache[2116];
endrule
rule s2118(sum_count == 2118);
  total_sum <= total_sum + cache[2117];
endrule
rule s2119(sum_count == 2119);
  total_sum <= total_sum + cache[2118];
endrule
rule s2120(sum_count == 2120);
  total_sum <= total_sum + cache[2119];
endrule
rule s2121(sum_count == 2121);
  total_sum <= total_sum + cache[2120];
endrule
rule s2122(sum_count == 2122);
  total_sum <= total_sum + cache[2121];
endrule
rule s2123(sum_count == 2123);
  total_sum <= total_sum + cache[2122];
endrule
rule s2124(sum_count == 2124);
  total_sum <= total_sum + cache[2123];
endrule
rule s2125(sum_count == 2125);
  total_sum <= total_sum + cache[2124];
endrule
rule s2126(sum_count == 2126);
  total_sum <= total_sum + cache[2125];
endrule
rule s2127(sum_count == 2127);
  total_sum <= total_sum + cache[2126];
endrule
rule s2128(sum_count == 2128);
  total_sum <= total_sum + cache[2127];
endrule
rule s2129(sum_count == 2129);
  total_sum <= total_sum + cache[2128];
endrule
rule s2130(sum_count == 2130);
  total_sum <= total_sum + cache[2129];
endrule
rule s2131(sum_count == 2131);
  total_sum <= total_sum + cache[2130];
endrule
rule s2132(sum_count == 2132);
  total_sum <= total_sum + cache[2131];
endrule
rule s2133(sum_count == 2133);
  total_sum <= total_sum + cache[2132];
endrule
rule s2134(sum_count == 2134);
  total_sum <= total_sum + cache[2133];
endrule
rule s2135(sum_count == 2135);
  total_sum <= total_sum + cache[2134];
endrule
rule s2136(sum_count == 2136);
  total_sum <= total_sum + cache[2135];
endrule
rule s2137(sum_count == 2137);
  total_sum <= total_sum + cache[2136];
endrule
rule s2138(sum_count == 2138);
  total_sum <= total_sum + cache[2137];
endrule
rule s2139(sum_count == 2139);
  total_sum <= total_sum + cache[2138];
endrule
rule s2140(sum_count == 2140);
  total_sum <= total_sum + cache[2139];
endrule
rule s2141(sum_count == 2141);
  total_sum <= total_sum + cache[2140];
endrule
rule s2142(sum_count == 2142);
  total_sum <= total_sum + cache[2141];
endrule
rule s2143(sum_count == 2143);
  total_sum <= total_sum + cache[2142];
endrule
rule s2144(sum_count == 2144);
  total_sum <= total_sum + cache[2143];
endrule
rule s2145(sum_count == 2145);
  total_sum <= total_sum + cache[2144];
endrule
rule s2146(sum_count == 2146);
  total_sum <= total_sum + cache[2145];
endrule
rule s2147(sum_count == 2147);
  total_sum <= total_sum + cache[2146];
endrule
rule s2148(sum_count == 2148);
  total_sum <= total_sum + cache[2147];
endrule
rule s2149(sum_count == 2149);
  total_sum <= total_sum + cache[2148];
endrule
rule s2150(sum_count == 2150);
  total_sum <= total_sum + cache[2149];
endrule
rule s2151(sum_count == 2151);
  total_sum <= total_sum + cache[2150];
endrule
rule s2152(sum_count == 2152);
  total_sum <= total_sum + cache[2151];
endrule
rule s2153(sum_count == 2153);
  total_sum <= total_sum + cache[2152];
endrule
rule s2154(sum_count == 2154);
  total_sum <= total_sum + cache[2153];
endrule
rule s2155(sum_count == 2155);
  total_sum <= total_sum + cache[2154];
endrule
rule s2156(sum_count == 2156);
  total_sum <= total_sum + cache[2155];
endrule
rule s2157(sum_count == 2157);
  total_sum <= total_sum + cache[2156];
endrule
rule s2158(sum_count == 2158);
  total_sum <= total_sum + cache[2157];
endrule
rule s2159(sum_count == 2159);
  total_sum <= total_sum + cache[2158];
endrule
rule s2160(sum_count == 2160);
  total_sum <= total_sum + cache[2159];
endrule
rule s2161(sum_count == 2161);
  total_sum <= total_sum + cache[2160];
endrule
rule s2162(sum_count == 2162);
  total_sum <= total_sum + cache[2161];
endrule
rule s2163(sum_count == 2163);
  total_sum <= total_sum + cache[2162];
endrule
rule s2164(sum_count == 2164);
  total_sum <= total_sum + cache[2163];
endrule
rule s2165(sum_count == 2165);
  total_sum <= total_sum + cache[2164];
endrule
rule s2166(sum_count == 2166);
  total_sum <= total_sum + cache[2165];
endrule
rule s2167(sum_count == 2167);
  total_sum <= total_sum + cache[2166];
endrule
rule s2168(sum_count == 2168);
  total_sum <= total_sum + cache[2167];
endrule
rule s2169(sum_count == 2169);
  total_sum <= total_sum + cache[2168];
endrule
rule s2170(sum_count == 2170);
  total_sum <= total_sum + cache[2169];
endrule
rule s2171(sum_count == 2171);
  total_sum <= total_sum + cache[2170];
endrule
rule s2172(sum_count == 2172);
  total_sum <= total_sum + cache[2171];
endrule
rule s2173(sum_count == 2173);
  total_sum <= total_sum + cache[2172];
endrule
rule s2174(sum_count == 2174);
  total_sum <= total_sum + cache[2173];
endrule
rule s2175(sum_count == 2175);
  total_sum <= total_sum + cache[2174];
endrule
rule s2176(sum_count == 2176);
  total_sum <= total_sum + cache[2175];
endrule
rule s2177(sum_count == 2177);
  total_sum <= total_sum + cache[2176];
endrule
rule s2178(sum_count == 2178);
  total_sum <= total_sum + cache[2177];
endrule
rule s2179(sum_count == 2179);
  total_sum <= total_sum + cache[2178];
endrule
rule s2180(sum_count == 2180);
  total_sum <= total_sum + cache[2179];
endrule
rule s2181(sum_count == 2181);
  total_sum <= total_sum + cache[2180];
endrule
rule s2182(sum_count == 2182);
  total_sum <= total_sum + cache[2181];
endrule
rule s2183(sum_count == 2183);
  total_sum <= total_sum + cache[2182];
endrule
rule s2184(sum_count == 2184);
  total_sum <= total_sum + cache[2183];
endrule
rule s2185(sum_count == 2185);
  total_sum <= total_sum + cache[2184];
endrule
rule s2186(sum_count == 2186);
  total_sum <= total_sum + cache[2185];
endrule
rule s2187(sum_count == 2187);
  total_sum <= total_sum + cache[2186];
endrule
rule s2188(sum_count == 2188);
  total_sum <= total_sum + cache[2187];
endrule
rule s2189(sum_count == 2189);
  total_sum <= total_sum + cache[2188];
endrule
rule s2190(sum_count == 2190);
  total_sum <= total_sum + cache[2189];
endrule
rule s2191(sum_count == 2191);
  total_sum <= total_sum + cache[2190];
endrule
rule s2192(sum_count == 2192);
  total_sum <= total_sum + cache[2191];
endrule
rule s2193(sum_count == 2193);
  total_sum <= total_sum + cache[2192];
endrule
rule s2194(sum_count == 2194);
  total_sum <= total_sum + cache[2193];
endrule
rule s2195(sum_count == 2195);
  total_sum <= total_sum + cache[2194];
endrule
rule s2196(sum_count == 2196);
  total_sum <= total_sum + cache[2195];
endrule
rule s2197(sum_count == 2197);
  total_sum <= total_sum + cache[2196];
endrule
rule s2198(sum_count == 2198);
  total_sum <= total_sum + cache[2197];
endrule
rule s2199(sum_count == 2199);
  total_sum <= total_sum + cache[2198];
endrule
rule s2200(sum_count == 2200);
  total_sum <= total_sum + cache[2199];
endrule
rule s2201(sum_count == 2201);
  total_sum <= total_sum + cache[2200];
endrule
rule s2202(sum_count == 2202);
  total_sum <= total_sum + cache[2201];
endrule
rule s2203(sum_count == 2203);
  total_sum <= total_sum + cache[2202];
endrule
rule s2204(sum_count == 2204);
  total_sum <= total_sum + cache[2203];
endrule
rule s2205(sum_count == 2205);
  total_sum <= total_sum + cache[2204];
endrule
rule s2206(sum_count == 2206);
  total_sum <= total_sum + cache[2205];
endrule
rule s2207(sum_count == 2207);
  total_sum <= total_sum + cache[2206];
endrule
rule s2208(sum_count == 2208);
  total_sum <= total_sum + cache[2207];
endrule
rule s2209(sum_count == 2209);
  total_sum <= total_sum + cache[2208];
endrule
rule s2210(sum_count == 2210);
  total_sum <= total_sum + cache[2209];
endrule
rule s2211(sum_count == 2211);
  total_sum <= total_sum + cache[2210];
endrule
rule s2212(sum_count == 2212);
  total_sum <= total_sum + cache[2211];
endrule
rule s2213(sum_count == 2213);
  total_sum <= total_sum + cache[2212];
endrule
rule s2214(sum_count == 2214);
  total_sum <= total_sum + cache[2213];
endrule
rule s2215(sum_count == 2215);
  total_sum <= total_sum + cache[2214];
endrule
rule s2216(sum_count == 2216);
  total_sum <= total_sum + cache[2215];
endrule
rule s2217(sum_count == 2217);
  total_sum <= total_sum + cache[2216];
endrule
rule s2218(sum_count == 2218);
  total_sum <= total_sum + cache[2217];
endrule
rule s2219(sum_count == 2219);
  total_sum <= total_sum + cache[2218];
endrule
rule s2220(sum_count == 2220);
  total_sum <= total_sum + cache[2219];
endrule
rule s2221(sum_count == 2221);
  total_sum <= total_sum + cache[2220];
endrule
rule s2222(sum_count == 2222);
  total_sum <= total_sum + cache[2221];
endrule
rule s2223(sum_count == 2223);
  total_sum <= total_sum + cache[2222];
endrule
rule s2224(sum_count == 2224);
  total_sum <= total_sum + cache[2223];
endrule
rule s2225(sum_count == 2225);
  total_sum <= total_sum + cache[2224];
endrule
rule s2226(sum_count == 2226);
  total_sum <= total_sum + cache[2225];
endrule
rule s2227(sum_count == 2227);
  total_sum <= total_sum + cache[2226];
endrule
rule s2228(sum_count == 2228);
  total_sum <= total_sum + cache[2227];
endrule
rule s2229(sum_count == 2229);
  total_sum <= total_sum + cache[2228];
endrule
rule s2230(sum_count == 2230);
  total_sum <= total_sum + cache[2229];
endrule
rule s2231(sum_count == 2231);
  total_sum <= total_sum + cache[2230];
endrule
rule s2232(sum_count == 2232);
  total_sum <= total_sum + cache[2231];
endrule
rule s2233(sum_count == 2233);
  total_sum <= total_sum + cache[2232];
endrule
rule s2234(sum_count == 2234);
  total_sum <= total_sum + cache[2233];
endrule
rule s2235(sum_count == 2235);
  total_sum <= total_sum + cache[2234];
endrule
rule s2236(sum_count == 2236);
  total_sum <= total_sum + cache[2235];
endrule
rule s2237(sum_count == 2237);
  total_sum <= total_sum + cache[2236];
endrule
rule s2238(sum_count == 2238);
  total_sum <= total_sum + cache[2237];
endrule
rule s2239(sum_count == 2239);
  total_sum <= total_sum + cache[2238];
endrule
rule s2240(sum_count == 2240);
  total_sum <= total_sum + cache[2239];
endrule
rule s2241(sum_count == 2241);
  total_sum <= total_sum + cache[2240];
endrule
rule s2242(sum_count == 2242);
  total_sum <= total_sum + cache[2241];
endrule
rule s2243(sum_count == 2243);
  total_sum <= total_sum + cache[2242];
endrule
rule s2244(sum_count == 2244);
  total_sum <= total_sum + cache[2243];
endrule
rule s2245(sum_count == 2245);
  total_sum <= total_sum + cache[2244];
endrule
rule s2246(sum_count == 2246);
  total_sum <= total_sum + cache[2245];
endrule
rule s2247(sum_count == 2247);
  total_sum <= total_sum + cache[2246];
endrule
rule s2248(sum_count == 2248);
  total_sum <= total_sum + cache[2247];
endrule
rule s2249(sum_count == 2249);
  total_sum <= total_sum + cache[2248];
endrule
rule s2250(sum_count == 2250);
  total_sum <= total_sum + cache[2249];
endrule
rule s2251(sum_count == 2251);
  total_sum <= total_sum + cache[2250];
endrule
rule s2252(sum_count == 2252);
  total_sum <= total_sum + cache[2251];
endrule
rule s2253(sum_count == 2253);
  total_sum <= total_sum + cache[2252];
endrule
rule s2254(sum_count == 2254);
  total_sum <= total_sum + cache[2253];
endrule
rule s2255(sum_count == 2255);
  total_sum <= total_sum + cache[2254];
endrule
rule s2256(sum_count == 2256);
  total_sum <= total_sum + cache[2255];
endrule
rule s2257(sum_count == 2257);
  total_sum <= total_sum + cache[2256];
endrule
rule s2258(sum_count == 2258);
  total_sum <= total_sum + cache[2257];
endrule
rule s2259(sum_count == 2259);
  total_sum <= total_sum + cache[2258];
endrule
rule s2260(sum_count == 2260);
  total_sum <= total_sum + cache[2259];
endrule
rule s2261(sum_count == 2261);
  total_sum <= total_sum + cache[2260];
endrule
rule s2262(sum_count == 2262);
  total_sum <= total_sum + cache[2261];
endrule
rule s2263(sum_count == 2263);
  total_sum <= total_sum + cache[2262];
endrule
rule s2264(sum_count == 2264);
  total_sum <= total_sum + cache[2263];
endrule
rule s2265(sum_count == 2265);
  total_sum <= total_sum + cache[2264];
endrule
rule s2266(sum_count == 2266);
  total_sum <= total_sum + cache[2265];
endrule
rule s2267(sum_count == 2267);
  total_sum <= total_sum + cache[2266];
endrule
rule s2268(sum_count == 2268);
  total_sum <= total_sum + cache[2267];
endrule
rule s2269(sum_count == 2269);
  total_sum <= total_sum + cache[2268];
endrule
rule s2270(sum_count == 2270);
  total_sum <= total_sum + cache[2269];
endrule
rule s2271(sum_count == 2271);
  total_sum <= total_sum + cache[2270];
endrule
rule s2272(sum_count == 2272);
  total_sum <= total_sum + cache[2271];
endrule
rule s2273(sum_count == 2273);
  total_sum <= total_sum + cache[2272];
endrule
rule s2274(sum_count == 2274);
  total_sum <= total_sum + cache[2273];
endrule
rule s2275(sum_count == 2275);
  total_sum <= total_sum + cache[2274];
endrule
rule s2276(sum_count == 2276);
  total_sum <= total_sum + cache[2275];
endrule
rule s2277(sum_count == 2277);
  total_sum <= total_sum + cache[2276];
endrule
rule s2278(sum_count == 2278);
  total_sum <= total_sum + cache[2277];
endrule
rule s2279(sum_count == 2279);
  total_sum <= total_sum + cache[2278];
endrule
rule s2280(sum_count == 2280);
  total_sum <= total_sum + cache[2279];
endrule
rule s2281(sum_count == 2281);
  total_sum <= total_sum + cache[2280];
endrule
rule s2282(sum_count == 2282);
  total_sum <= total_sum + cache[2281];
endrule
rule s2283(sum_count == 2283);
  total_sum <= total_sum + cache[2282];
endrule
rule s2284(sum_count == 2284);
  total_sum <= total_sum + cache[2283];
endrule
rule s2285(sum_count == 2285);
  total_sum <= total_sum + cache[2284];
endrule
rule s2286(sum_count == 2286);
  total_sum <= total_sum + cache[2285];
endrule
rule s2287(sum_count == 2287);
  total_sum <= total_sum + cache[2286];
endrule
rule s2288(sum_count == 2288);
  total_sum <= total_sum + cache[2287];
endrule
rule s2289(sum_count == 2289);
  total_sum <= total_sum + cache[2288];
endrule
rule s2290(sum_count == 2290);
  total_sum <= total_sum + cache[2289];
endrule
rule s2291(sum_count == 2291);
  total_sum <= total_sum + cache[2290];
endrule
rule s2292(sum_count == 2292);
  total_sum <= total_sum + cache[2291];
endrule
rule s2293(sum_count == 2293);
  total_sum <= total_sum + cache[2292];
endrule
rule s2294(sum_count == 2294);
  total_sum <= total_sum + cache[2293];
endrule
rule s2295(sum_count == 2295);
  total_sum <= total_sum + cache[2294];
endrule
rule s2296(sum_count == 2296);
  total_sum <= total_sum + cache[2295];
endrule
rule s2297(sum_count == 2297);
  total_sum <= total_sum + cache[2296];
endrule
rule s2298(sum_count == 2298);
  total_sum <= total_sum + cache[2297];
endrule
rule s2299(sum_count == 2299);
  total_sum <= total_sum + cache[2298];
endrule
rule s2300(sum_count == 2300);
  total_sum <= total_sum + cache[2299];
endrule
rule s2301(sum_count == 2301);
  total_sum <= total_sum + cache[2300];
endrule
rule s2302(sum_count == 2302);
  total_sum <= total_sum + cache[2301];
endrule
rule s2303(sum_count == 2303);
  total_sum <= total_sum + cache[2302];
endrule
rule s2304(sum_count == 2304);
  total_sum <= total_sum + cache[2303];
endrule
rule s2305(sum_count == 2305);
  total_sum <= total_sum + cache[2304];
endrule
rule s2306(sum_count == 2306);
  total_sum <= total_sum + cache[2305];
endrule
rule s2307(sum_count == 2307);
  total_sum <= total_sum + cache[2306];
endrule
rule s2308(sum_count == 2308);
  total_sum <= total_sum + cache[2307];
endrule
rule s2309(sum_count == 2309);
  total_sum <= total_sum + cache[2308];
endrule
rule s2310(sum_count == 2310);
  total_sum <= total_sum + cache[2309];
endrule
rule s2311(sum_count == 2311);
  total_sum <= total_sum + cache[2310];
endrule
rule s2312(sum_count == 2312);
  total_sum <= total_sum + cache[2311];
endrule
rule s2313(sum_count == 2313);
  total_sum <= total_sum + cache[2312];
endrule
rule s2314(sum_count == 2314);
  total_sum <= total_sum + cache[2313];
endrule
rule s2315(sum_count == 2315);
  total_sum <= total_sum + cache[2314];
endrule
rule s2316(sum_count == 2316);
  total_sum <= total_sum + cache[2315];
endrule
rule s2317(sum_count == 2317);
  total_sum <= total_sum + cache[2316];
endrule
rule s2318(sum_count == 2318);
  total_sum <= total_sum + cache[2317];
endrule
rule s2319(sum_count == 2319);
  total_sum <= total_sum + cache[2318];
endrule
rule s2320(sum_count == 2320);
  total_sum <= total_sum + cache[2319];
endrule
rule s2321(sum_count == 2321);
  total_sum <= total_sum + cache[2320];
endrule
rule s2322(sum_count == 2322);
  total_sum <= total_sum + cache[2321];
endrule
rule s2323(sum_count == 2323);
  total_sum <= total_sum + cache[2322];
endrule
rule s2324(sum_count == 2324);
  total_sum <= total_sum + cache[2323];
endrule
rule s2325(sum_count == 2325);
  total_sum <= total_sum + cache[2324];
endrule
rule s2326(sum_count == 2326);
  total_sum <= total_sum + cache[2325];
endrule
rule s2327(sum_count == 2327);
  total_sum <= total_sum + cache[2326];
endrule
rule s2328(sum_count == 2328);
  total_sum <= total_sum + cache[2327];
endrule
rule s2329(sum_count == 2329);
  total_sum <= total_sum + cache[2328];
endrule
rule s2330(sum_count == 2330);
  total_sum <= total_sum + cache[2329];
endrule
rule s2331(sum_count == 2331);
  total_sum <= total_sum + cache[2330];
endrule
rule s2332(sum_count == 2332);
  total_sum <= total_sum + cache[2331];
endrule
rule s2333(sum_count == 2333);
  total_sum <= total_sum + cache[2332];
endrule
rule s2334(sum_count == 2334);
  total_sum <= total_sum + cache[2333];
endrule
rule s2335(sum_count == 2335);
  total_sum <= total_sum + cache[2334];
endrule
rule s2336(sum_count == 2336);
  total_sum <= total_sum + cache[2335];
endrule
rule s2337(sum_count == 2337);
  total_sum <= total_sum + cache[2336];
endrule
rule s2338(sum_count == 2338);
  total_sum <= total_sum + cache[2337];
endrule
rule s2339(sum_count == 2339);
  total_sum <= total_sum + cache[2338];
endrule
rule s2340(sum_count == 2340);
  total_sum <= total_sum + cache[2339];
endrule
rule s2341(sum_count == 2341);
  total_sum <= total_sum + cache[2340];
endrule
rule s2342(sum_count == 2342);
  total_sum <= total_sum + cache[2341];
endrule
rule s2343(sum_count == 2343);
  total_sum <= total_sum + cache[2342];
endrule
rule s2344(sum_count == 2344);
  total_sum <= total_sum + cache[2343];
endrule
rule s2345(sum_count == 2345);
  total_sum <= total_sum + cache[2344];
endrule
rule s2346(sum_count == 2346);
  total_sum <= total_sum + cache[2345];
endrule
rule s2347(sum_count == 2347);
  total_sum <= total_sum + cache[2346];
endrule
rule s2348(sum_count == 2348);
  total_sum <= total_sum + cache[2347];
endrule
rule s2349(sum_count == 2349);
  total_sum <= total_sum + cache[2348];
endrule
rule s2350(sum_count == 2350);
  total_sum <= total_sum + cache[2349];
endrule
rule s2351(sum_count == 2351);
  total_sum <= total_sum + cache[2350];
endrule
rule s2352(sum_count == 2352);
  total_sum <= total_sum + cache[2351];
endrule
rule s2353(sum_count == 2353);
  total_sum <= total_sum + cache[2352];
endrule
rule s2354(sum_count == 2354);
  total_sum <= total_sum + cache[2353];
endrule
rule s2355(sum_count == 2355);
  total_sum <= total_sum + cache[2354];
endrule
rule s2356(sum_count == 2356);
  total_sum <= total_sum + cache[2355];
endrule
rule s2357(sum_count == 2357);
  total_sum <= total_sum + cache[2356];
endrule
rule s2358(sum_count == 2358);
  total_sum <= total_sum + cache[2357];
endrule
rule s2359(sum_count == 2359);
  total_sum <= total_sum + cache[2358];
endrule
rule s2360(sum_count == 2360);
  total_sum <= total_sum + cache[2359];
endrule
rule s2361(sum_count == 2361);
  total_sum <= total_sum + cache[2360];
endrule
rule s2362(sum_count == 2362);
  total_sum <= total_sum + cache[2361];
endrule
rule s2363(sum_count == 2363);
  total_sum <= total_sum + cache[2362];
endrule
rule s2364(sum_count == 2364);
  total_sum <= total_sum + cache[2363];
endrule
rule s2365(sum_count == 2365);
  total_sum <= total_sum + cache[2364];
endrule
rule s2366(sum_count == 2366);
  total_sum <= total_sum + cache[2365];
endrule
rule s2367(sum_count == 2367);
  total_sum <= total_sum + cache[2366];
endrule
rule s2368(sum_count == 2368);
  total_sum <= total_sum + cache[2367];
endrule
rule s2369(sum_count == 2369);
  total_sum <= total_sum + cache[2368];
endrule
rule s2370(sum_count == 2370);
  total_sum <= total_sum + cache[2369];
endrule
rule s2371(sum_count == 2371);
  total_sum <= total_sum + cache[2370];
endrule
rule s2372(sum_count == 2372);
  total_sum <= total_sum + cache[2371];
endrule
rule s2373(sum_count == 2373);
  total_sum <= total_sum + cache[2372];
endrule
rule s2374(sum_count == 2374);
  total_sum <= total_sum + cache[2373];
endrule
rule s2375(sum_count == 2375);
  total_sum <= total_sum + cache[2374];
endrule
rule s2376(sum_count == 2376);
  total_sum <= total_sum + cache[2375];
endrule
rule s2377(sum_count == 2377);
  total_sum <= total_sum + cache[2376];
endrule
rule s2378(sum_count == 2378);
  total_sum <= total_sum + cache[2377];
endrule
rule s2379(sum_count == 2379);
  total_sum <= total_sum + cache[2378];
endrule
rule s2380(sum_count == 2380);
  total_sum <= total_sum + cache[2379];
endrule
rule s2381(sum_count == 2381);
  total_sum <= total_sum + cache[2380];
endrule
rule s2382(sum_count == 2382);
  total_sum <= total_sum + cache[2381];
endrule
rule s2383(sum_count == 2383);
  total_sum <= total_sum + cache[2382];
endrule
rule s2384(sum_count == 2384);
  total_sum <= total_sum + cache[2383];
endrule
rule s2385(sum_count == 2385);
  total_sum <= total_sum + cache[2384];
endrule
rule s2386(sum_count == 2386);
  total_sum <= total_sum + cache[2385];
endrule
rule s2387(sum_count == 2387);
  total_sum <= total_sum + cache[2386];
endrule
rule s2388(sum_count == 2388);
  total_sum <= total_sum + cache[2387];
endrule
rule s2389(sum_count == 2389);
  total_sum <= total_sum + cache[2388];
endrule
rule s2390(sum_count == 2390);
  total_sum <= total_sum + cache[2389];
endrule
rule s2391(sum_count == 2391);
  total_sum <= total_sum + cache[2390];
endrule
rule s2392(sum_count == 2392);
  total_sum <= total_sum + cache[2391];
endrule
rule s2393(sum_count == 2393);
  total_sum <= total_sum + cache[2392];
endrule
rule s2394(sum_count == 2394);
  total_sum <= total_sum + cache[2393];
endrule
rule s2395(sum_count == 2395);
  total_sum <= total_sum + cache[2394];
endrule
rule s2396(sum_count == 2396);
  total_sum <= total_sum + cache[2395];
endrule
rule s2397(sum_count == 2397);
  total_sum <= total_sum + cache[2396];
endrule
rule s2398(sum_count == 2398);
  total_sum <= total_sum + cache[2397];
endrule
rule s2399(sum_count == 2399);
  total_sum <= total_sum + cache[2398];
endrule
rule s2400(sum_count == 2400);
  total_sum <= total_sum + cache[2399];
endrule
rule s2401(sum_count == 2401);
  total_sum <= total_sum + cache[2400];
endrule
rule s2402(sum_count == 2402);
  total_sum <= total_sum + cache[2401];
endrule
rule s2403(sum_count == 2403);
  total_sum <= total_sum + cache[2402];
endrule
rule s2404(sum_count == 2404);
  total_sum <= total_sum + cache[2403];
endrule
rule s2405(sum_count == 2405);
  total_sum <= total_sum + cache[2404];
endrule
rule s2406(sum_count == 2406);
  total_sum <= total_sum + cache[2405];
endrule
rule s2407(sum_count == 2407);
  total_sum <= total_sum + cache[2406];
endrule
rule s2408(sum_count == 2408);
  total_sum <= total_sum + cache[2407];
endrule
rule s2409(sum_count == 2409);
  total_sum <= total_sum + cache[2408];
endrule
rule s2410(sum_count == 2410);
  total_sum <= total_sum + cache[2409];
endrule
rule s2411(sum_count == 2411);
  total_sum <= total_sum + cache[2410];
endrule
rule s2412(sum_count == 2412);
  total_sum <= total_sum + cache[2411];
endrule
rule s2413(sum_count == 2413);
  total_sum <= total_sum + cache[2412];
endrule
rule s2414(sum_count == 2414);
  total_sum <= total_sum + cache[2413];
endrule
rule s2415(sum_count == 2415);
  total_sum <= total_sum + cache[2414];
endrule
rule s2416(sum_count == 2416);
  total_sum <= total_sum + cache[2415];
endrule
rule s2417(sum_count == 2417);
  total_sum <= total_sum + cache[2416];
endrule
rule s2418(sum_count == 2418);
  total_sum <= total_sum + cache[2417];
endrule
rule s2419(sum_count == 2419);
  total_sum <= total_sum + cache[2418];
endrule
rule s2420(sum_count == 2420);
  total_sum <= total_sum + cache[2419];
endrule
rule s2421(sum_count == 2421);
  total_sum <= total_sum + cache[2420];
endrule
rule s2422(sum_count == 2422);
  total_sum <= total_sum + cache[2421];
endrule
rule s2423(sum_count == 2423);
  total_sum <= total_sum + cache[2422];
endrule
rule s2424(sum_count == 2424);
  total_sum <= total_sum + cache[2423];
endrule
rule s2425(sum_count == 2425);
  total_sum <= total_sum + cache[2424];
endrule
rule s2426(sum_count == 2426);
  total_sum <= total_sum + cache[2425];
endrule
rule s2427(sum_count == 2427);
  total_sum <= total_sum + cache[2426];
endrule
rule s2428(sum_count == 2428);
  total_sum <= total_sum + cache[2427];
endrule
rule s2429(sum_count == 2429);
  total_sum <= total_sum + cache[2428];
endrule
rule s2430(sum_count == 2430);
  total_sum <= total_sum + cache[2429];
endrule
rule s2431(sum_count == 2431);
  total_sum <= total_sum + cache[2430];
endrule
rule s2432(sum_count == 2432);
  total_sum <= total_sum + cache[2431];
endrule
rule s2433(sum_count == 2433);
  total_sum <= total_sum + cache[2432];
endrule
rule s2434(sum_count == 2434);
  total_sum <= total_sum + cache[2433];
endrule
rule s2435(sum_count == 2435);
  total_sum <= total_sum + cache[2434];
endrule
rule s2436(sum_count == 2436);
  total_sum <= total_sum + cache[2435];
endrule
rule s2437(sum_count == 2437);
  total_sum <= total_sum + cache[2436];
endrule
rule s2438(sum_count == 2438);
  total_sum <= total_sum + cache[2437];
endrule
rule s2439(sum_count == 2439);
  total_sum <= total_sum + cache[2438];
endrule
rule s2440(sum_count == 2440);
  total_sum <= total_sum + cache[2439];
endrule
rule s2441(sum_count == 2441);
  total_sum <= total_sum + cache[2440];
endrule
rule s2442(sum_count == 2442);
  total_sum <= total_sum + cache[2441];
endrule
rule s2443(sum_count == 2443);
  total_sum <= total_sum + cache[2442];
endrule
rule s2444(sum_count == 2444);
  total_sum <= total_sum + cache[2443];
endrule
rule s2445(sum_count == 2445);
  total_sum <= total_sum + cache[2444];
endrule
rule s2446(sum_count == 2446);
  total_sum <= total_sum + cache[2445];
endrule
rule s2447(sum_count == 2447);
  total_sum <= total_sum + cache[2446];
endrule
rule s2448(sum_count == 2448);
  total_sum <= total_sum + cache[2447];
endrule
rule s2449(sum_count == 2449);
  total_sum <= total_sum + cache[2448];
endrule
rule s2450(sum_count == 2450);
  total_sum <= total_sum + cache[2449];
endrule
rule s2451(sum_count == 2451);
  total_sum <= total_sum + cache[2450];
endrule
rule s2452(sum_count == 2452);
  total_sum <= total_sum + cache[2451];
endrule
rule s2453(sum_count == 2453);
  total_sum <= total_sum + cache[2452];
endrule
rule s2454(sum_count == 2454);
  total_sum <= total_sum + cache[2453];
endrule
rule s2455(sum_count == 2455);
  total_sum <= total_sum + cache[2454];
endrule
rule s2456(sum_count == 2456);
  total_sum <= total_sum + cache[2455];
endrule
rule s2457(sum_count == 2457);
  total_sum <= total_sum + cache[2456];
endrule
rule s2458(sum_count == 2458);
  total_sum <= total_sum + cache[2457];
endrule
rule s2459(sum_count == 2459);
  total_sum <= total_sum + cache[2458];
endrule
rule s2460(sum_count == 2460);
  total_sum <= total_sum + cache[2459];
endrule
rule s2461(sum_count == 2461);
  total_sum <= total_sum + cache[2460];
endrule
rule s2462(sum_count == 2462);
  total_sum <= total_sum + cache[2461];
endrule
rule s2463(sum_count == 2463);
  total_sum <= total_sum + cache[2462];
endrule
rule s2464(sum_count == 2464);
  total_sum <= total_sum + cache[2463];
endrule
rule s2465(sum_count == 2465);
  total_sum <= total_sum + cache[2464];
endrule
rule s2466(sum_count == 2466);
  total_sum <= total_sum + cache[2465];
endrule
rule s2467(sum_count == 2467);
  total_sum <= total_sum + cache[2466];
endrule
rule s2468(sum_count == 2468);
  total_sum <= total_sum + cache[2467];
endrule
rule s2469(sum_count == 2469);
  total_sum <= total_sum + cache[2468];
endrule
rule s2470(sum_count == 2470);
  total_sum <= total_sum + cache[2469];
endrule
rule s2471(sum_count == 2471);
  total_sum <= total_sum + cache[2470];
endrule
rule s2472(sum_count == 2472);
  total_sum <= total_sum + cache[2471];
endrule
rule s2473(sum_count == 2473);
  total_sum <= total_sum + cache[2472];
endrule
rule s2474(sum_count == 2474);
  total_sum <= total_sum + cache[2473];
endrule
rule s2475(sum_count == 2475);
  total_sum <= total_sum + cache[2474];
endrule
rule s2476(sum_count == 2476);
  total_sum <= total_sum + cache[2475];
endrule
rule s2477(sum_count == 2477);
  total_sum <= total_sum + cache[2476];
endrule
rule s2478(sum_count == 2478);
  total_sum <= total_sum + cache[2477];
endrule
rule s2479(sum_count == 2479);
  total_sum <= total_sum + cache[2478];
endrule
rule s2480(sum_count == 2480);
  total_sum <= total_sum + cache[2479];
endrule
rule s2481(sum_count == 2481);
  total_sum <= total_sum + cache[2480];
endrule
rule s2482(sum_count == 2482);
  total_sum <= total_sum + cache[2481];
endrule
rule s2483(sum_count == 2483);
  total_sum <= total_sum + cache[2482];
endrule
rule s2484(sum_count == 2484);
  total_sum <= total_sum + cache[2483];
endrule
rule s2485(sum_count == 2485);
  total_sum <= total_sum + cache[2484];
endrule
rule s2486(sum_count == 2486);
  total_sum <= total_sum + cache[2485];
endrule
rule s2487(sum_count == 2487);
  total_sum <= total_sum + cache[2486];
endrule
rule s2488(sum_count == 2488);
  total_sum <= total_sum + cache[2487];
endrule
rule s2489(sum_count == 2489);
  total_sum <= total_sum + cache[2488];
endrule
rule s2490(sum_count == 2490);
  total_sum <= total_sum + cache[2489];
endrule
rule s2491(sum_count == 2491);
  total_sum <= total_sum + cache[2490];
endrule
rule s2492(sum_count == 2492);
  total_sum <= total_sum + cache[2491];
endrule
rule s2493(sum_count == 2493);
  total_sum <= total_sum + cache[2492];
endrule
rule s2494(sum_count == 2494);
  total_sum <= total_sum + cache[2493];
endrule
rule s2495(sum_count == 2495);
  total_sum <= total_sum + cache[2494];
endrule
rule s2496(sum_count == 2496);
  total_sum <= total_sum + cache[2495];
endrule
rule s2497(sum_count == 2497);
  total_sum <= total_sum + cache[2496];
endrule
rule s2498(sum_count == 2498);
  total_sum <= total_sum + cache[2497];
endrule
rule s2499(sum_count == 2499);
  total_sum <= total_sum + cache[2498];
endrule
rule s2500(sum_count == 2500);
  total_sum <= total_sum + cache[2499];
endrule
rule s2501(sum_count == 2501);
  total_sum <= total_sum + cache[2500];
endrule
rule s2502(sum_count == 2502);
  total_sum <= total_sum + cache[2501];
endrule
rule s2503(sum_count == 2503);
  total_sum <= total_sum + cache[2502];
endrule
rule s2504(sum_count == 2504);
  total_sum <= total_sum + cache[2503];
endrule
rule s2505(sum_count == 2505);
  total_sum <= total_sum + cache[2504];
endrule
rule s2506(sum_count == 2506);
  total_sum <= total_sum + cache[2505];
endrule
rule s2507(sum_count == 2507);
  total_sum <= total_sum + cache[2506];
endrule
rule s2508(sum_count == 2508);
  total_sum <= total_sum + cache[2507];
endrule
rule s2509(sum_count == 2509);
  total_sum <= total_sum + cache[2508];
endrule
rule s2510(sum_count == 2510);
  total_sum <= total_sum + cache[2509];
endrule
rule s2511(sum_count == 2511);
  total_sum <= total_sum + cache[2510];
endrule
rule s2512(sum_count == 2512);
  total_sum <= total_sum + cache[2511];
endrule
rule s2513(sum_count == 2513);
  total_sum <= total_sum + cache[2512];
endrule
rule s2514(sum_count == 2514);
  total_sum <= total_sum + cache[2513];
endrule
rule s2515(sum_count == 2515);
  total_sum <= total_sum + cache[2514];
endrule
rule s2516(sum_count == 2516);
  total_sum <= total_sum + cache[2515];
endrule
rule s2517(sum_count == 2517);
  total_sum <= total_sum + cache[2516];
endrule
rule s2518(sum_count == 2518);
  total_sum <= total_sum + cache[2517];
endrule
rule s2519(sum_count == 2519);
  total_sum <= total_sum + cache[2518];
endrule
rule s2520(sum_count == 2520);
  total_sum <= total_sum + cache[2519];
endrule
rule s2521(sum_count == 2521);
  total_sum <= total_sum + cache[2520];
endrule
rule s2522(sum_count == 2522);
  total_sum <= total_sum + cache[2521];
endrule
rule s2523(sum_count == 2523);
  total_sum <= total_sum + cache[2522];
endrule
rule s2524(sum_count == 2524);
  total_sum <= total_sum + cache[2523];
endrule
rule s2525(sum_count == 2525);
  total_sum <= total_sum + cache[2524];
endrule
rule s2526(sum_count == 2526);
  total_sum <= total_sum + cache[2525];
endrule
rule s2527(sum_count == 2527);
  total_sum <= total_sum + cache[2526];
endrule
rule s2528(sum_count == 2528);
  total_sum <= total_sum + cache[2527];
endrule
rule s2529(sum_count == 2529);
  total_sum <= total_sum + cache[2528];
endrule
rule s2530(sum_count == 2530);
  total_sum <= total_sum + cache[2529];
endrule
rule s2531(sum_count == 2531);
  total_sum <= total_sum + cache[2530];
endrule
rule s2532(sum_count == 2532);
  total_sum <= total_sum + cache[2531];
endrule
rule s2533(sum_count == 2533);
  total_sum <= total_sum + cache[2532];
endrule
rule s2534(sum_count == 2534);
  total_sum <= total_sum + cache[2533];
endrule
rule s2535(sum_count == 2535);
  total_sum <= total_sum + cache[2534];
endrule
rule s2536(sum_count == 2536);
  total_sum <= total_sum + cache[2535];
endrule
rule s2537(sum_count == 2537);
  total_sum <= total_sum + cache[2536];
endrule
rule s2538(sum_count == 2538);
  total_sum <= total_sum + cache[2537];
endrule
rule s2539(sum_count == 2539);
  total_sum <= total_sum + cache[2538];
endrule
rule s2540(sum_count == 2540);
  total_sum <= total_sum + cache[2539];
endrule
rule s2541(sum_count == 2541);
  total_sum <= total_sum + cache[2540];
endrule
rule s2542(sum_count == 2542);
  total_sum <= total_sum + cache[2541];
endrule
rule s2543(sum_count == 2543);
  total_sum <= total_sum + cache[2542];
endrule
rule s2544(sum_count == 2544);
  total_sum <= total_sum + cache[2543];
endrule
rule s2545(sum_count == 2545);
  total_sum <= total_sum + cache[2544];
endrule
rule s2546(sum_count == 2546);
  total_sum <= total_sum + cache[2545];
endrule
rule s2547(sum_count == 2547);
  total_sum <= total_sum + cache[2546];
endrule
rule s2548(sum_count == 2548);
  total_sum <= total_sum + cache[2547];
endrule
rule s2549(sum_count == 2549);
  total_sum <= total_sum + cache[2548];
endrule
rule s2550(sum_count == 2550);
  total_sum <= total_sum + cache[2549];
endrule
rule s2551(sum_count == 2551);
  total_sum <= total_sum + cache[2550];
endrule
rule s2552(sum_count == 2552);
  total_sum <= total_sum + cache[2551];
endrule
rule s2553(sum_count == 2553);
  total_sum <= total_sum + cache[2552];
endrule
rule s2554(sum_count == 2554);
  total_sum <= total_sum + cache[2553];
endrule
rule s2555(sum_count == 2555);
  total_sum <= total_sum + cache[2554];
endrule
rule s2556(sum_count == 2556);
  total_sum <= total_sum + cache[2555];
endrule
rule s2557(sum_count == 2557);
  total_sum <= total_sum + cache[2556];
endrule
rule s2558(sum_count == 2558);
  total_sum <= total_sum + cache[2557];
endrule
rule s2559(sum_count == 2559);
  total_sum <= total_sum + cache[2558];
endrule
rule s2560(sum_count == 2560);
  total_sum <= total_sum + cache[2559];
endrule
rule s2561(sum_count == 2561);
  total_sum <= total_sum + cache[2560];
endrule
rule s2562(sum_count == 2562);
  total_sum <= total_sum + cache[2561];
endrule
rule s2563(sum_count == 2563);
  total_sum <= total_sum + cache[2562];
endrule
rule s2564(sum_count == 2564);
  total_sum <= total_sum + cache[2563];
endrule
rule s2565(sum_count == 2565);
  total_sum <= total_sum + cache[2564];
endrule
rule s2566(sum_count == 2566);
  total_sum <= total_sum + cache[2565];
endrule
rule s2567(sum_count == 2567);
  total_sum <= total_sum + cache[2566];
endrule
rule s2568(sum_count == 2568);
  total_sum <= total_sum + cache[2567];
endrule
rule s2569(sum_count == 2569);
  total_sum <= total_sum + cache[2568];
endrule
rule s2570(sum_count == 2570);
  total_sum <= total_sum + cache[2569];
endrule
rule s2571(sum_count == 2571);
  total_sum <= total_sum + cache[2570];
endrule
rule s2572(sum_count == 2572);
  total_sum <= total_sum + cache[2571];
endrule
rule s2573(sum_count == 2573);
  total_sum <= total_sum + cache[2572];
endrule
rule s2574(sum_count == 2574);
  total_sum <= total_sum + cache[2573];
endrule
rule s2575(sum_count == 2575);
  total_sum <= total_sum + cache[2574];
endrule
rule s2576(sum_count == 2576);
  total_sum <= total_sum + cache[2575];
endrule
rule s2577(sum_count == 2577);
  total_sum <= total_sum + cache[2576];
endrule
rule s2578(sum_count == 2578);
  total_sum <= total_sum + cache[2577];
endrule
rule s2579(sum_count == 2579);
  total_sum <= total_sum + cache[2578];
endrule
rule s2580(sum_count == 2580);
  total_sum <= total_sum + cache[2579];
endrule
rule s2581(sum_count == 2581);
  total_sum <= total_sum + cache[2580];
endrule
rule s2582(sum_count == 2582);
  total_sum <= total_sum + cache[2581];
endrule
rule s2583(sum_count == 2583);
  total_sum <= total_sum + cache[2582];
endrule
rule s2584(sum_count == 2584);
  total_sum <= total_sum + cache[2583];
endrule
rule s2585(sum_count == 2585);
  total_sum <= total_sum + cache[2584];
endrule
rule s2586(sum_count == 2586);
  total_sum <= total_sum + cache[2585];
endrule
rule s2587(sum_count == 2587);
  total_sum <= total_sum + cache[2586];
endrule
rule s2588(sum_count == 2588);
  total_sum <= total_sum + cache[2587];
endrule
rule s2589(sum_count == 2589);
  total_sum <= total_sum + cache[2588];
endrule
rule s2590(sum_count == 2590);
  total_sum <= total_sum + cache[2589];
endrule
rule s2591(sum_count == 2591);
  total_sum <= total_sum + cache[2590];
endrule
rule s2592(sum_count == 2592);
  total_sum <= total_sum + cache[2591];
endrule
rule s2593(sum_count == 2593);
  total_sum <= total_sum + cache[2592];
endrule
rule s2594(sum_count == 2594);
  total_sum <= total_sum + cache[2593];
endrule
rule s2595(sum_count == 2595);
  total_sum <= total_sum + cache[2594];
endrule
rule s2596(sum_count == 2596);
  total_sum <= total_sum + cache[2595];
endrule
rule s2597(sum_count == 2597);
  total_sum <= total_sum + cache[2596];
endrule
rule s2598(sum_count == 2598);
  total_sum <= total_sum + cache[2597];
endrule
rule s2599(sum_count == 2599);
  total_sum <= total_sum + cache[2598];
endrule
rule s2600(sum_count == 2600);
  total_sum <= total_sum + cache[2599];
endrule
rule s2601(sum_count == 2601);
  total_sum <= total_sum + cache[2600];
endrule
rule s2602(sum_count == 2602);
  total_sum <= total_sum + cache[2601];
endrule
rule s2603(sum_count == 2603);
  total_sum <= total_sum + cache[2602];
endrule
rule s2604(sum_count == 2604);
  total_sum <= total_sum + cache[2603];
endrule
rule s2605(sum_count == 2605);
  total_sum <= total_sum + cache[2604];
endrule
rule s2606(sum_count == 2606);
  total_sum <= total_sum + cache[2605];
endrule
rule s2607(sum_count == 2607);
  total_sum <= total_sum + cache[2606];
endrule
rule s2608(sum_count == 2608);
  total_sum <= total_sum + cache[2607];
endrule
rule s2609(sum_count == 2609);
  total_sum <= total_sum + cache[2608];
endrule
rule s2610(sum_count == 2610);
  total_sum <= total_sum + cache[2609];
endrule
rule s2611(sum_count == 2611);
  total_sum <= total_sum + cache[2610];
endrule
rule s2612(sum_count == 2612);
  total_sum <= total_sum + cache[2611];
endrule
rule s2613(sum_count == 2613);
  total_sum <= total_sum + cache[2612];
endrule
rule s2614(sum_count == 2614);
  total_sum <= total_sum + cache[2613];
endrule
rule s2615(sum_count == 2615);
  total_sum <= total_sum + cache[2614];
endrule
rule s2616(sum_count == 2616);
  total_sum <= total_sum + cache[2615];
endrule
rule s2617(sum_count == 2617);
  total_sum <= total_sum + cache[2616];
endrule
rule s2618(sum_count == 2618);
  total_sum <= total_sum + cache[2617];
endrule
rule s2619(sum_count == 2619);
  total_sum <= total_sum + cache[2618];
endrule
rule s2620(sum_count == 2620);
  total_sum <= total_sum + cache[2619];
endrule
rule s2621(sum_count == 2621);
  total_sum <= total_sum + cache[2620];
endrule
rule s2622(sum_count == 2622);
  total_sum <= total_sum + cache[2621];
endrule
rule s2623(sum_count == 2623);
  total_sum <= total_sum + cache[2622];
endrule
rule s2624(sum_count == 2624);
  total_sum <= total_sum + cache[2623];
endrule
rule s2625(sum_count == 2625);
  total_sum <= total_sum + cache[2624];
endrule
rule s2626(sum_count == 2626);
  total_sum <= total_sum + cache[2625];
endrule
rule s2627(sum_count == 2627);
  total_sum <= total_sum + cache[2626];
endrule
rule s2628(sum_count == 2628);
  total_sum <= total_sum + cache[2627];
endrule
rule s2629(sum_count == 2629);
  total_sum <= total_sum + cache[2628];
endrule
rule s2630(sum_count == 2630);
  total_sum <= total_sum + cache[2629];
endrule
rule s2631(sum_count == 2631);
  total_sum <= total_sum + cache[2630];
endrule
rule s2632(sum_count == 2632);
  total_sum <= total_sum + cache[2631];
endrule
rule s2633(sum_count == 2633);
  total_sum <= total_sum + cache[2632];
endrule
rule s2634(sum_count == 2634);
  total_sum <= total_sum + cache[2633];
endrule
rule s2635(sum_count == 2635);
  total_sum <= total_sum + cache[2634];
endrule
rule s2636(sum_count == 2636);
  total_sum <= total_sum + cache[2635];
endrule
rule s2637(sum_count == 2637);
  total_sum <= total_sum + cache[2636];
endrule
rule s2638(sum_count == 2638);
  total_sum <= total_sum + cache[2637];
endrule
rule s2639(sum_count == 2639);
  total_sum <= total_sum + cache[2638];
endrule
rule s2640(sum_count == 2640);
  total_sum <= total_sum + cache[2639];
endrule
rule s2641(sum_count == 2641);
  total_sum <= total_sum + cache[2640];
endrule
rule s2642(sum_count == 2642);
  total_sum <= total_sum + cache[2641];
endrule
rule s2643(sum_count == 2643);
  total_sum <= total_sum + cache[2642];
endrule
rule s2644(sum_count == 2644);
  total_sum <= total_sum + cache[2643];
endrule
rule s2645(sum_count == 2645);
  total_sum <= total_sum + cache[2644];
endrule
rule s2646(sum_count == 2646);
  total_sum <= total_sum + cache[2645];
endrule
rule s2647(sum_count == 2647);
  total_sum <= total_sum + cache[2646];
endrule
rule s2648(sum_count == 2648);
  total_sum <= total_sum + cache[2647];
endrule
rule s2649(sum_count == 2649);
  total_sum <= total_sum + cache[2648];
endrule
rule s2650(sum_count == 2650);
  total_sum <= total_sum + cache[2649];
endrule
rule s2651(sum_count == 2651);
  total_sum <= total_sum + cache[2650];
endrule
rule s2652(sum_count == 2652);
  total_sum <= total_sum + cache[2651];
endrule
rule s2653(sum_count == 2653);
  total_sum <= total_sum + cache[2652];
endrule
rule s2654(sum_count == 2654);
  total_sum <= total_sum + cache[2653];
endrule
rule s2655(sum_count == 2655);
  total_sum <= total_sum + cache[2654];
endrule
rule s2656(sum_count == 2656);
  total_sum <= total_sum + cache[2655];
endrule
rule s2657(sum_count == 2657);
  total_sum <= total_sum + cache[2656];
endrule
rule s2658(sum_count == 2658);
  total_sum <= total_sum + cache[2657];
endrule
rule s2659(sum_count == 2659);
  total_sum <= total_sum + cache[2658];
endrule
rule s2660(sum_count == 2660);
  total_sum <= total_sum + cache[2659];
endrule
rule s2661(sum_count == 2661);
  total_sum <= total_sum + cache[2660];
endrule
rule s2662(sum_count == 2662);
  total_sum <= total_sum + cache[2661];
endrule
rule s2663(sum_count == 2663);
  total_sum <= total_sum + cache[2662];
endrule
rule s2664(sum_count == 2664);
  total_sum <= total_sum + cache[2663];
endrule
rule s2665(sum_count == 2665);
  total_sum <= total_sum + cache[2664];
endrule
rule s2666(sum_count == 2666);
  total_sum <= total_sum + cache[2665];
endrule
rule s2667(sum_count == 2667);
  total_sum <= total_sum + cache[2666];
endrule
rule s2668(sum_count == 2668);
  total_sum <= total_sum + cache[2667];
endrule
rule s2669(sum_count == 2669);
  total_sum <= total_sum + cache[2668];
endrule
rule s2670(sum_count == 2670);
  total_sum <= total_sum + cache[2669];
endrule
rule s2671(sum_count == 2671);
  total_sum <= total_sum + cache[2670];
endrule
rule s2672(sum_count == 2672);
  total_sum <= total_sum + cache[2671];
endrule
rule s2673(sum_count == 2673);
  total_sum <= total_sum + cache[2672];
endrule
rule s2674(sum_count == 2674);
  total_sum <= total_sum + cache[2673];
endrule
rule s2675(sum_count == 2675);
  total_sum <= total_sum + cache[2674];
endrule
rule s2676(sum_count == 2676);
  total_sum <= total_sum + cache[2675];
endrule
rule s2677(sum_count == 2677);
  total_sum <= total_sum + cache[2676];
endrule
rule s2678(sum_count == 2678);
  total_sum <= total_sum + cache[2677];
endrule
rule s2679(sum_count == 2679);
  total_sum <= total_sum + cache[2678];
endrule
rule s2680(sum_count == 2680);
  total_sum <= total_sum + cache[2679];
endrule
rule s2681(sum_count == 2681);
  total_sum <= total_sum + cache[2680];
endrule
rule s2682(sum_count == 2682);
  total_sum <= total_sum + cache[2681];
endrule
rule s2683(sum_count == 2683);
  total_sum <= total_sum + cache[2682];
endrule
rule s2684(sum_count == 2684);
  total_sum <= total_sum + cache[2683];
endrule
rule s2685(sum_count == 2685);
  total_sum <= total_sum + cache[2684];
endrule
rule s2686(sum_count == 2686);
  total_sum <= total_sum + cache[2685];
endrule
rule s2687(sum_count == 2687);
  total_sum <= total_sum + cache[2686];
endrule
rule s2688(sum_count == 2688);
  total_sum <= total_sum + cache[2687];
endrule
rule s2689(sum_count == 2689);
  total_sum <= total_sum + cache[2688];
endrule
rule s2690(sum_count == 2690);
  total_sum <= total_sum + cache[2689];
endrule
rule s2691(sum_count == 2691);
  total_sum <= total_sum + cache[2690];
endrule
rule s2692(sum_count == 2692);
  total_sum <= total_sum + cache[2691];
endrule
rule s2693(sum_count == 2693);
  total_sum <= total_sum + cache[2692];
endrule
rule s2694(sum_count == 2694);
  total_sum <= total_sum + cache[2693];
endrule
rule s2695(sum_count == 2695);
  total_sum <= total_sum + cache[2694];
endrule
rule s2696(sum_count == 2696);
  total_sum <= total_sum + cache[2695];
endrule
rule s2697(sum_count == 2697);
  total_sum <= total_sum + cache[2696];
endrule
rule s2698(sum_count == 2698);
  total_sum <= total_sum + cache[2697];
endrule
rule s2699(sum_count == 2699);
  total_sum <= total_sum + cache[2698];
endrule
rule s2700(sum_count == 2700);
  total_sum <= total_sum + cache[2699];
endrule
rule s2701(sum_count == 2701);
  total_sum <= total_sum + cache[2700];
endrule
rule s2702(sum_count == 2702);
  total_sum <= total_sum + cache[2701];
endrule
rule s2703(sum_count == 2703);
  total_sum <= total_sum + cache[2702];
endrule
rule s2704(sum_count == 2704);
  total_sum <= total_sum + cache[2703];
endrule
rule s2705(sum_count == 2705);
  total_sum <= total_sum + cache[2704];
endrule
rule s2706(sum_count == 2706);
  total_sum <= total_sum + cache[2705];
endrule
rule s2707(sum_count == 2707);
  total_sum <= total_sum + cache[2706];
endrule
rule s2708(sum_count == 2708);
  total_sum <= total_sum + cache[2707];
endrule
rule s2709(sum_count == 2709);
  total_sum <= total_sum + cache[2708];
endrule
rule s2710(sum_count == 2710);
  total_sum <= total_sum + cache[2709];
endrule
rule s2711(sum_count == 2711);
  total_sum <= total_sum + cache[2710];
endrule
rule s2712(sum_count == 2712);
  total_sum <= total_sum + cache[2711];
endrule
rule s2713(sum_count == 2713);
  total_sum <= total_sum + cache[2712];
endrule
rule s2714(sum_count == 2714);
  total_sum <= total_sum + cache[2713];
endrule
rule s2715(sum_count == 2715);
  total_sum <= total_sum + cache[2714];
endrule
rule s2716(sum_count == 2716);
  total_sum <= total_sum + cache[2715];
endrule
rule s2717(sum_count == 2717);
  total_sum <= total_sum + cache[2716];
endrule
rule s2718(sum_count == 2718);
  total_sum <= total_sum + cache[2717];
endrule
rule s2719(sum_count == 2719);
  total_sum <= total_sum + cache[2718];
endrule
rule s2720(sum_count == 2720);
  total_sum <= total_sum + cache[2719];
endrule
rule s2721(sum_count == 2721);
  total_sum <= total_sum + cache[2720];
endrule
rule s2722(sum_count == 2722);
  total_sum <= total_sum + cache[2721];
endrule
rule s2723(sum_count == 2723);
  total_sum <= total_sum + cache[2722];
endrule
rule s2724(sum_count == 2724);
  total_sum <= total_sum + cache[2723];
endrule
rule s2725(sum_count == 2725);
  total_sum <= total_sum + cache[2724];
endrule
rule s2726(sum_count == 2726);
  total_sum <= total_sum + cache[2725];
endrule
rule s2727(sum_count == 2727);
  total_sum <= total_sum + cache[2726];
endrule
rule s2728(sum_count == 2728);
  total_sum <= total_sum + cache[2727];
endrule
rule s2729(sum_count == 2729);
  total_sum <= total_sum + cache[2728];
endrule
rule s2730(sum_count == 2730);
  total_sum <= total_sum + cache[2729];
endrule
rule s2731(sum_count == 2731);
  total_sum <= total_sum + cache[2730];
endrule
rule s2732(sum_count == 2732);
  total_sum <= total_sum + cache[2731];
endrule
rule s2733(sum_count == 2733);
  total_sum <= total_sum + cache[2732];
endrule
rule s2734(sum_count == 2734);
  total_sum <= total_sum + cache[2733];
endrule
rule s2735(sum_count == 2735);
  total_sum <= total_sum + cache[2734];
endrule
rule s2736(sum_count == 2736);
  total_sum <= total_sum + cache[2735];
endrule
rule s2737(sum_count == 2737);
  total_sum <= total_sum + cache[2736];
endrule
rule s2738(sum_count == 2738);
  total_sum <= total_sum + cache[2737];
endrule
rule s2739(sum_count == 2739);
  total_sum <= total_sum + cache[2738];
endrule
rule s2740(sum_count == 2740);
  total_sum <= total_sum + cache[2739];
endrule
rule s2741(sum_count == 2741);
  total_sum <= total_sum + cache[2740];
endrule
rule s2742(sum_count == 2742);
  total_sum <= total_sum + cache[2741];
endrule
rule s2743(sum_count == 2743);
  total_sum <= total_sum + cache[2742];
endrule
rule s2744(sum_count == 2744);
  total_sum <= total_sum + cache[2743];
endrule
rule s2745(sum_count == 2745);
  total_sum <= total_sum + cache[2744];
endrule
rule s2746(sum_count == 2746);
  total_sum <= total_sum + cache[2745];
endrule
rule s2747(sum_count == 2747);
  total_sum <= total_sum + cache[2746];
endrule
rule s2748(sum_count == 2748);
  total_sum <= total_sum + cache[2747];
endrule
rule s2749(sum_count == 2749);
  total_sum <= total_sum + cache[2748];
endrule
rule s2750(sum_count == 2750);
  total_sum <= total_sum + cache[2749];
endrule
rule s2751(sum_count == 2751);
  total_sum <= total_sum + cache[2750];
endrule
rule s2752(sum_count == 2752);
  total_sum <= total_sum + cache[2751];
endrule
rule s2753(sum_count == 2753);
  total_sum <= total_sum + cache[2752];
endrule
rule s2754(sum_count == 2754);
  total_sum <= total_sum + cache[2753];
endrule
rule s2755(sum_count == 2755);
  total_sum <= total_sum + cache[2754];
endrule
rule s2756(sum_count == 2756);
  total_sum <= total_sum + cache[2755];
endrule
rule s2757(sum_count == 2757);
  total_sum <= total_sum + cache[2756];
endrule
rule s2758(sum_count == 2758);
  total_sum <= total_sum + cache[2757];
endrule
rule s2759(sum_count == 2759);
  total_sum <= total_sum + cache[2758];
endrule
rule s2760(sum_count == 2760);
  total_sum <= total_sum + cache[2759];
endrule
rule s2761(sum_count == 2761);
  total_sum <= total_sum + cache[2760];
endrule
rule s2762(sum_count == 2762);
  total_sum <= total_sum + cache[2761];
endrule
rule s2763(sum_count == 2763);
  total_sum <= total_sum + cache[2762];
endrule
rule s2764(sum_count == 2764);
  total_sum <= total_sum + cache[2763];
endrule
rule s2765(sum_count == 2765);
  total_sum <= total_sum + cache[2764];
endrule
rule s2766(sum_count == 2766);
  total_sum <= total_sum + cache[2765];
endrule
rule s2767(sum_count == 2767);
  total_sum <= total_sum + cache[2766];
endrule
rule s2768(sum_count == 2768);
  total_sum <= total_sum + cache[2767];
endrule
rule s2769(sum_count == 2769);
  total_sum <= total_sum + cache[2768];
endrule
rule s2770(sum_count == 2770);
  total_sum <= total_sum + cache[2769];
endrule
rule s2771(sum_count == 2771);
  total_sum <= total_sum + cache[2770];
endrule
rule s2772(sum_count == 2772);
  total_sum <= total_sum + cache[2771];
endrule
rule s2773(sum_count == 2773);
  total_sum <= total_sum + cache[2772];
endrule
rule s2774(sum_count == 2774);
  total_sum <= total_sum + cache[2773];
endrule
rule s2775(sum_count == 2775);
  total_sum <= total_sum + cache[2774];
endrule
rule s2776(sum_count == 2776);
  total_sum <= total_sum + cache[2775];
endrule
rule s2777(sum_count == 2777);
  total_sum <= total_sum + cache[2776];
endrule
rule s2778(sum_count == 2778);
  total_sum <= total_sum + cache[2777];
endrule
rule s2779(sum_count == 2779);
  total_sum <= total_sum + cache[2778];
endrule
rule s2780(sum_count == 2780);
  total_sum <= total_sum + cache[2779];
endrule
rule s2781(sum_count == 2781);
  total_sum <= total_sum + cache[2780];
endrule
rule s2782(sum_count == 2782);
  total_sum <= total_sum + cache[2781];
endrule
rule s2783(sum_count == 2783);
  total_sum <= total_sum + cache[2782];
endrule
rule s2784(sum_count == 2784);
  total_sum <= total_sum + cache[2783];
endrule
rule s2785(sum_count == 2785);
  total_sum <= total_sum + cache[2784];
endrule
rule s2786(sum_count == 2786);
  total_sum <= total_sum + cache[2785];
endrule
rule s2787(sum_count == 2787);
  total_sum <= total_sum + cache[2786];
endrule
rule s2788(sum_count == 2788);
  total_sum <= total_sum + cache[2787];
endrule
rule s2789(sum_count == 2789);
  total_sum <= total_sum + cache[2788];
endrule
rule s2790(sum_count == 2790);
  total_sum <= total_sum + cache[2789];
endrule
rule s2791(sum_count == 2791);
  total_sum <= total_sum + cache[2790];
endrule
rule s2792(sum_count == 2792);
  total_sum <= total_sum + cache[2791];
endrule
rule s2793(sum_count == 2793);
  total_sum <= total_sum + cache[2792];
endrule
rule s2794(sum_count == 2794);
  total_sum <= total_sum + cache[2793];
endrule
rule s2795(sum_count == 2795);
  total_sum <= total_sum + cache[2794];
endrule
rule s2796(sum_count == 2796);
  total_sum <= total_sum + cache[2795];
endrule
rule s2797(sum_count == 2797);
  total_sum <= total_sum + cache[2796];
endrule
rule s2798(sum_count == 2798);
  total_sum <= total_sum + cache[2797];
endrule
rule s2799(sum_count == 2799);
  total_sum <= total_sum + cache[2798];
endrule
rule s2800(sum_count == 2800);
  total_sum <= total_sum + cache[2799];
endrule
rule s2801(sum_count == 2801);
  total_sum <= total_sum + cache[2800];
endrule
rule s2802(sum_count == 2802);
  total_sum <= total_sum + cache[2801];
endrule
rule s2803(sum_count == 2803);
  total_sum <= total_sum + cache[2802];
endrule
rule s2804(sum_count == 2804);
  total_sum <= total_sum + cache[2803];
endrule
rule s2805(sum_count == 2805);
  total_sum <= total_sum + cache[2804];
endrule
rule s2806(sum_count == 2806);
  total_sum <= total_sum + cache[2805];
endrule
rule s2807(sum_count == 2807);
  total_sum <= total_sum + cache[2806];
endrule
rule s2808(sum_count == 2808);
  total_sum <= total_sum + cache[2807];
endrule
rule s2809(sum_count == 2809);
  total_sum <= total_sum + cache[2808];
endrule
rule s2810(sum_count == 2810);
  total_sum <= total_sum + cache[2809];
endrule
rule s2811(sum_count == 2811);
  total_sum <= total_sum + cache[2810];
endrule
rule s2812(sum_count == 2812);
  total_sum <= total_sum + cache[2811];
endrule
rule s2813(sum_count == 2813);
  total_sum <= total_sum + cache[2812];
endrule
rule s2814(sum_count == 2814);
  total_sum <= total_sum + cache[2813];
endrule
rule s2815(sum_count == 2815);
  total_sum <= total_sum + cache[2814];
endrule
rule s2816(sum_count == 2816);
  total_sum <= total_sum + cache[2815];
endrule
rule s2817(sum_count == 2817);
  total_sum <= total_sum + cache[2816];
endrule
rule s2818(sum_count == 2818);
  total_sum <= total_sum + cache[2817];
endrule
rule s2819(sum_count == 2819);
  total_sum <= total_sum + cache[2818];
endrule
rule s2820(sum_count == 2820);
  total_sum <= total_sum + cache[2819];
endrule
rule s2821(sum_count == 2821);
  total_sum <= total_sum + cache[2820];
endrule
rule s2822(sum_count == 2822);
  total_sum <= total_sum + cache[2821];
endrule
rule s2823(sum_count == 2823);
  total_sum <= total_sum + cache[2822];
endrule
rule s2824(sum_count == 2824);
  total_sum <= total_sum + cache[2823];
endrule
rule s2825(sum_count == 2825);
  total_sum <= total_sum + cache[2824];
endrule
rule s2826(sum_count == 2826);
  total_sum <= total_sum + cache[2825];
endrule
rule s2827(sum_count == 2827);
  total_sum <= total_sum + cache[2826];
endrule
rule s2828(sum_count == 2828);
  total_sum <= total_sum + cache[2827];
endrule
rule s2829(sum_count == 2829);
  total_sum <= total_sum + cache[2828];
endrule
rule s2830(sum_count == 2830);
  total_sum <= total_sum + cache[2829];
endrule
rule s2831(sum_count == 2831);
  total_sum <= total_sum + cache[2830];
endrule
rule s2832(sum_count == 2832);
  total_sum <= total_sum + cache[2831];
endrule
rule s2833(sum_count == 2833);
  total_sum <= total_sum + cache[2832];
endrule
rule s2834(sum_count == 2834);
  total_sum <= total_sum + cache[2833];
endrule
rule s2835(sum_count == 2835);
  total_sum <= total_sum + cache[2834];
endrule
rule s2836(sum_count == 2836);
  total_sum <= total_sum + cache[2835];
endrule
rule s2837(sum_count == 2837);
  total_sum <= total_sum + cache[2836];
endrule
rule s2838(sum_count == 2838);
  total_sum <= total_sum + cache[2837];
endrule
rule s2839(sum_count == 2839);
  total_sum <= total_sum + cache[2838];
endrule
rule s2840(sum_count == 2840);
  total_sum <= total_sum + cache[2839];
endrule
rule s2841(sum_count == 2841);
  total_sum <= total_sum + cache[2840];
endrule
rule s2842(sum_count == 2842);
  total_sum <= total_sum + cache[2841];
endrule
rule s2843(sum_count == 2843);
  total_sum <= total_sum + cache[2842];
endrule
rule s2844(sum_count == 2844);
  total_sum <= total_sum + cache[2843];
endrule
rule s2845(sum_count == 2845);
  total_sum <= total_sum + cache[2844];
endrule
rule s2846(sum_count == 2846);
  total_sum <= total_sum + cache[2845];
endrule
rule s2847(sum_count == 2847);
  total_sum <= total_sum + cache[2846];
endrule
rule s2848(sum_count == 2848);
  total_sum <= total_sum + cache[2847];
endrule
rule s2849(sum_count == 2849);
  total_sum <= total_sum + cache[2848];
endrule
rule s2850(sum_count == 2850);
  total_sum <= total_sum + cache[2849];
endrule
rule s2851(sum_count == 2851);
  total_sum <= total_sum + cache[2850];
endrule
rule s2852(sum_count == 2852);
  total_sum <= total_sum + cache[2851];
endrule
rule s2853(sum_count == 2853);
  total_sum <= total_sum + cache[2852];
endrule
rule s2854(sum_count == 2854);
  total_sum <= total_sum + cache[2853];
endrule
rule s2855(sum_count == 2855);
  total_sum <= total_sum + cache[2854];
endrule
rule s2856(sum_count == 2856);
  total_sum <= total_sum + cache[2855];
endrule
rule s2857(sum_count == 2857);
  total_sum <= total_sum + cache[2856];
endrule
rule s2858(sum_count == 2858);
  total_sum <= total_sum + cache[2857];
endrule
rule s2859(sum_count == 2859);
  total_sum <= total_sum + cache[2858];
endrule
rule s2860(sum_count == 2860);
  total_sum <= total_sum + cache[2859];
endrule
rule s2861(sum_count == 2861);
  total_sum <= total_sum + cache[2860];
endrule
rule s2862(sum_count == 2862);
  total_sum <= total_sum + cache[2861];
endrule
rule s2863(sum_count == 2863);
  total_sum <= total_sum + cache[2862];
endrule
rule s2864(sum_count == 2864);
  total_sum <= total_sum + cache[2863];
endrule
rule s2865(sum_count == 2865);
  total_sum <= total_sum + cache[2864];
endrule
rule s2866(sum_count == 2866);
  total_sum <= total_sum + cache[2865];
endrule
rule s2867(sum_count == 2867);
  total_sum <= total_sum + cache[2866];
endrule
rule s2868(sum_count == 2868);
  total_sum <= total_sum + cache[2867];
endrule
rule s2869(sum_count == 2869);
  total_sum <= total_sum + cache[2868];
endrule
rule s2870(sum_count == 2870);
  total_sum <= total_sum + cache[2869];
endrule
rule s2871(sum_count == 2871);
  total_sum <= total_sum + cache[2870];
endrule
rule s2872(sum_count == 2872);
  total_sum <= total_sum + cache[2871];
endrule
rule s2873(sum_count == 2873);
  total_sum <= total_sum + cache[2872];
endrule
rule s2874(sum_count == 2874);
  total_sum <= total_sum + cache[2873];
endrule
rule s2875(sum_count == 2875);
  total_sum <= total_sum + cache[2874];
endrule
rule s2876(sum_count == 2876);
  total_sum <= total_sum + cache[2875];
endrule
rule s2877(sum_count == 2877);
  total_sum <= total_sum + cache[2876];
endrule
rule s2878(sum_count == 2878);
  total_sum <= total_sum + cache[2877];
endrule
rule s2879(sum_count == 2879);
  total_sum <= total_sum + cache[2878];
endrule
rule s2880(sum_count == 2880);
  total_sum <= total_sum + cache[2879];
endrule
rule s2881(sum_count == 2881);
  total_sum <= total_sum + cache[2880];
endrule
rule s2882(sum_count == 2882);
  total_sum <= total_sum + cache[2881];
endrule
rule s2883(sum_count == 2883);
  total_sum <= total_sum + cache[2882];
endrule
rule s2884(sum_count == 2884);
  total_sum <= total_sum + cache[2883];
endrule
rule s2885(sum_count == 2885);
  total_sum <= total_sum + cache[2884];
endrule
rule s2886(sum_count == 2886);
  total_sum <= total_sum + cache[2885];
endrule
rule s2887(sum_count == 2887);
  total_sum <= total_sum + cache[2886];
endrule
rule s2888(sum_count == 2888);
  total_sum <= total_sum + cache[2887];
endrule
rule s2889(sum_count == 2889);
  total_sum <= total_sum + cache[2888];
endrule
rule s2890(sum_count == 2890);
  total_sum <= total_sum + cache[2889];
endrule
rule s2891(sum_count == 2891);
  total_sum <= total_sum + cache[2890];
endrule
rule s2892(sum_count == 2892);
  total_sum <= total_sum + cache[2891];
endrule
rule s2893(sum_count == 2893);
  total_sum <= total_sum + cache[2892];
endrule
rule s2894(sum_count == 2894);
  total_sum <= total_sum + cache[2893];
endrule
rule s2895(sum_count == 2895);
  total_sum <= total_sum + cache[2894];
endrule
rule s2896(sum_count == 2896);
  total_sum <= total_sum + cache[2895];
endrule
rule s2897(sum_count == 2897);
  total_sum <= total_sum + cache[2896];
endrule
rule s2898(sum_count == 2898);
  total_sum <= total_sum + cache[2897];
endrule
rule s2899(sum_count == 2899);
  total_sum <= total_sum + cache[2898];
endrule
rule s2900(sum_count == 2900);
  total_sum <= total_sum + cache[2899];
endrule
rule s2901(sum_count == 2901);
  total_sum <= total_sum + cache[2900];
endrule
rule s2902(sum_count == 2902);
  total_sum <= total_sum + cache[2901];
endrule
rule s2903(sum_count == 2903);
  total_sum <= total_sum + cache[2902];
endrule
rule s2904(sum_count == 2904);
  total_sum <= total_sum + cache[2903];
endrule
rule s2905(sum_count == 2905);
  total_sum <= total_sum + cache[2904];
endrule
rule s2906(sum_count == 2906);
  total_sum <= total_sum + cache[2905];
endrule
rule s2907(sum_count == 2907);
  total_sum <= total_sum + cache[2906];
endrule
rule s2908(sum_count == 2908);
  total_sum <= total_sum + cache[2907];
endrule
rule s2909(sum_count == 2909);
  total_sum <= total_sum + cache[2908];
endrule
rule s2910(sum_count == 2910);
  total_sum <= total_sum + cache[2909];
endrule
rule s2911(sum_count == 2911);
  total_sum <= total_sum + cache[2910];
endrule
rule s2912(sum_count == 2912);
  total_sum <= total_sum + cache[2911];
endrule
rule s2913(sum_count == 2913);
  total_sum <= total_sum + cache[2912];
endrule
rule s2914(sum_count == 2914);
  total_sum <= total_sum + cache[2913];
endrule
rule s2915(sum_count == 2915);
  total_sum <= total_sum + cache[2914];
endrule
rule s2916(sum_count == 2916);
  total_sum <= total_sum + cache[2915];
endrule
rule s2917(sum_count == 2917);
  total_sum <= total_sum + cache[2916];
endrule
rule s2918(sum_count == 2918);
  total_sum <= total_sum + cache[2917];
endrule
rule s2919(sum_count == 2919);
  total_sum <= total_sum + cache[2918];
endrule
rule s2920(sum_count == 2920);
  total_sum <= total_sum + cache[2919];
endrule
rule s2921(sum_count == 2921);
  total_sum <= total_sum + cache[2920];
endrule
rule s2922(sum_count == 2922);
  total_sum <= total_sum + cache[2921];
endrule
rule s2923(sum_count == 2923);
  total_sum <= total_sum + cache[2922];
endrule
rule s2924(sum_count == 2924);
  total_sum <= total_sum + cache[2923];
endrule
rule s2925(sum_count == 2925);
  total_sum <= total_sum + cache[2924];
endrule
rule s2926(sum_count == 2926);
  total_sum <= total_sum + cache[2925];
endrule
rule s2927(sum_count == 2927);
  total_sum <= total_sum + cache[2926];
endrule
rule s2928(sum_count == 2928);
  total_sum <= total_sum + cache[2927];
endrule
rule s2929(sum_count == 2929);
  total_sum <= total_sum + cache[2928];
endrule
rule s2930(sum_count == 2930);
  total_sum <= total_sum + cache[2929];
endrule
rule s2931(sum_count == 2931);
  total_sum <= total_sum + cache[2930];
endrule
rule s2932(sum_count == 2932);
  total_sum <= total_sum + cache[2931];
endrule
rule s2933(sum_count == 2933);
  total_sum <= total_sum + cache[2932];
endrule
rule s2934(sum_count == 2934);
  total_sum <= total_sum + cache[2933];
endrule
rule s2935(sum_count == 2935);
  total_sum <= total_sum + cache[2934];
endrule
rule s2936(sum_count == 2936);
  total_sum <= total_sum + cache[2935];
endrule
rule s2937(sum_count == 2937);
  total_sum <= total_sum + cache[2936];
endrule
rule s2938(sum_count == 2938);
  total_sum <= total_sum + cache[2937];
endrule
rule s2939(sum_count == 2939);
  total_sum <= total_sum + cache[2938];
endrule
rule s2940(sum_count == 2940);
  total_sum <= total_sum + cache[2939];
endrule
rule s2941(sum_count == 2941);
  total_sum <= total_sum + cache[2940];
endrule
rule s2942(sum_count == 2942);
  total_sum <= total_sum + cache[2941];
endrule
rule s2943(sum_count == 2943);
  total_sum <= total_sum + cache[2942];
endrule
rule s2944(sum_count == 2944);
  total_sum <= total_sum + cache[2943];
endrule
rule s2945(sum_count == 2945);
  total_sum <= total_sum + cache[2944];
endrule
rule s2946(sum_count == 2946);
  total_sum <= total_sum + cache[2945];
endrule
rule s2947(sum_count == 2947);
  total_sum <= total_sum + cache[2946];
endrule
rule s2948(sum_count == 2948);
  total_sum <= total_sum + cache[2947];
endrule
rule s2949(sum_count == 2949);
  total_sum <= total_sum + cache[2948];
endrule
rule s2950(sum_count == 2950);
  total_sum <= total_sum + cache[2949];
endrule
rule s2951(sum_count == 2951);
  total_sum <= total_sum + cache[2950];
endrule
rule s2952(sum_count == 2952);
  total_sum <= total_sum + cache[2951];
endrule
rule s2953(sum_count == 2953);
  total_sum <= total_sum + cache[2952];
endrule
rule s2954(sum_count == 2954);
  total_sum <= total_sum + cache[2953];
endrule
rule s2955(sum_count == 2955);
  total_sum <= total_sum + cache[2954];
endrule
rule s2956(sum_count == 2956);
  total_sum <= total_sum + cache[2955];
endrule
rule s2957(sum_count == 2957);
  total_sum <= total_sum + cache[2956];
endrule
rule s2958(sum_count == 2958);
  total_sum <= total_sum + cache[2957];
endrule
rule s2959(sum_count == 2959);
  total_sum <= total_sum + cache[2958];
endrule
rule s2960(sum_count == 2960);
  total_sum <= total_sum + cache[2959];
endrule
rule s2961(sum_count == 2961);
  total_sum <= total_sum + cache[2960];
endrule
rule s2962(sum_count == 2962);
  total_sum <= total_sum + cache[2961];
endrule
rule s2963(sum_count == 2963);
  total_sum <= total_sum + cache[2962];
endrule
rule s2964(sum_count == 2964);
  total_sum <= total_sum + cache[2963];
endrule
rule s2965(sum_count == 2965);
  total_sum <= total_sum + cache[2964];
endrule
rule s2966(sum_count == 2966);
  total_sum <= total_sum + cache[2965];
endrule
rule s2967(sum_count == 2967);
  total_sum <= total_sum + cache[2966];
endrule
rule s2968(sum_count == 2968);
  total_sum <= total_sum + cache[2967];
endrule
rule s2969(sum_count == 2969);
  total_sum <= total_sum + cache[2968];
endrule
rule s2970(sum_count == 2970);
  total_sum <= total_sum + cache[2969];
endrule
rule s2971(sum_count == 2971);
  total_sum <= total_sum + cache[2970];
endrule
rule s2972(sum_count == 2972);
  total_sum <= total_sum + cache[2971];
endrule
rule s2973(sum_count == 2973);
  total_sum <= total_sum + cache[2972];
endrule
rule s2974(sum_count == 2974);
  total_sum <= total_sum + cache[2973];
endrule
rule s2975(sum_count == 2975);
  total_sum <= total_sum + cache[2974];
endrule
rule s2976(sum_count == 2976);
  total_sum <= total_sum + cache[2975];
endrule
rule s2977(sum_count == 2977);
  total_sum <= total_sum + cache[2976];
endrule
rule s2978(sum_count == 2978);
  total_sum <= total_sum + cache[2977];
endrule
rule s2979(sum_count == 2979);
  total_sum <= total_sum + cache[2978];
endrule
rule s2980(sum_count == 2980);
  total_sum <= total_sum + cache[2979];
endrule
rule s2981(sum_count == 2981);
  total_sum <= total_sum + cache[2980];
endrule
rule s2982(sum_count == 2982);
  total_sum <= total_sum + cache[2981];
endrule
rule s2983(sum_count == 2983);
  total_sum <= total_sum + cache[2982];
endrule
rule s2984(sum_count == 2984);
  total_sum <= total_sum + cache[2983];
endrule
rule s2985(sum_count == 2985);
  total_sum <= total_sum + cache[2984];
endrule
rule s2986(sum_count == 2986);
  total_sum <= total_sum + cache[2985];
endrule
rule s2987(sum_count == 2987);
  total_sum <= total_sum + cache[2986];
endrule
rule s2988(sum_count == 2988);
  total_sum <= total_sum + cache[2987];
endrule
rule s2989(sum_count == 2989);
  total_sum <= total_sum + cache[2988];
endrule
rule s2990(sum_count == 2990);
  total_sum <= total_sum + cache[2989];
endrule
rule s2991(sum_count == 2991);
  total_sum <= total_sum + cache[2990];
endrule
rule s2992(sum_count == 2992);
  total_sum <= total_sum + cache[2991];
endrule
rule s2993(sum_count == 2993);
  total_sum <= total_sum + cache[2992];
endrule
rule s2994(sum_count == 2994);
  total_sum <= total_sum + cache[2993];
endrule
rule s2995(sum_count == 2995);
  total_sum <= total_sum + cache[2994];
endrule
rule s2996(sum_count == 2996);
  total_sum <= total_sum + cache[2995];
endrule
rule s2997(sum_count == 2997);
  total_sum <= total_sum + cache[2996];
endrule
rule s2998(sum_count == 2998);
  total_sum <= total_sum + cache[2997];
endrule
rule s2999(sum_count == 2999);
  total_sum <= total_sum + cache[2998];
endrule
rule s3000(sum_count == 3000);
  total_sum <= total_sum + cache[2999];
endrule
rule s3001(sum_count == 3001);
  total_sum <= total_sum + cache[3000];
endrule
rule s3002(sum_count == 3002);
  total_sum <= total_sum + cache[3001];
endrule
rule s3003(sum_count == 3003);
  total_sum <= total_sum + cache[3002];
endrule
rule s3004(sum_count == 3004);
  total_sum <= total_sum + cache[3003];
endrule
rule s3005(sum_count == 3005);
  total_sum <= total_sum + cache[3004];
endrule
rule s3006(sum_count == 3006);
  total_sum <= total_sum + cache[3005];
endrule
rule s3007(sum_count == 3007);
  total_sum <= total_sum + cache[3006];
endrule
rule s3008(sum_count == 3008);
  total_sum <= total_sum + cache[3007];
endrule
rule s3009(sum_count == 3009);
  total_sum <= total_sum + cache[3008];
endrule
rule s3010(sum_count == 3010);
  total_sum <= total_sum + cache[3009];
endrule
rule s3011(sum_count == 3011);
  total_sum <= total_sum + cache[3010];
endrule
rule s3012(sum_count == 3012);
  total_sum <= total_sum + cache[3011];
endrule
rule s3013(sum_count == 3013);
  total_sum <= total_sum + cache[3012];
endrule
rule s3014(sum_count == 3014);
  total_sum <= total_sum + cache[3013];
endrule
rule s3015(sum_count == 3015);
  total_sum <= total_sum + cache[3014];
endrule
rule s3016(sum_count == 3016);
  total_sum <= total_sum + cache[3015];
endrule
rule s3017(sum_count == 3017);
  total_sum <= total_sum + cache[3016];
endrule
rule s3018(sum_count == 3018);
  total_sum <= total_sum + cache[3017];
endrule
rule s3019(sum_count == 3019);
  total_sum <= total_sum + cache[3018];
endrule
rule s3020(sum_count == 3020);
  total_sum <= total_sum + cache[3019];
endrule
rule s3021(sum_count == 3021);
  total_sum <= total_sum + cache[3020];
endrule
rule s3022(sum_count == 3022);
  total_sum <= total_sum + cache[3021];
endrule
rule s3023(sum_count == 3023);
  total_sum <= total_sum + cache[3022];
endrule
rule s3024(sum_count == 3024);
  total_sum <= total_sum + cache[3023];
endrule
rule s3025(sum_count == 3025);
  total_sum <= total_sum + cache[3024];
endrule
rule s3026(sum_count == 3026);
  total_sum <= total_sum + cache[3025];
endrule
rule s3027(sum_count == 3027);
  total_sum <= total_sum + cache[3026];
endrule
rule s3028(sum_count == 3028);
  total_sum <= total_sum + cache[3027];
endrule
rule s3029(sum_count == 3029);
  total_sum <= total_sum + cache[3028];
endrule
rule s3030(sum_count == 3030);
  total_sum <= total_sum + cache[3029];
endrule
rule s3031(sum_count == 3031);
  total_sum <= total_sum + cache[3030];
endrule
rule s3032(sum_count == 3032);
  total_sum <= total_sum + cache[3031];
endrule
rule s3033(sum_count == 3033);
  total_sum <= total_sum + cache[3032];
endrule
rule s3034(sum_count == 3034);
  total_sum <= total_sum + cache[3033];
endrule
rule s3035(sum_count == 3035);
  total_sum <= total_sum + cache[3034];
endrule
rule s3036(sum_count == 3036);
  total_sum <= total_sum + cache[3035];
endrule
rule s3037(sum_count == 3037);
  total_sum <= total_sum + cache[3036];
endrule
rule s3038(sum_count == 3038);
  total_sum <= total_sum + cache[3037];
endrule
rule s3039(sum_count == 3039);
  total_sum <= total_sum + cache[3038];
endrule
rule s3040(sum_count == 3040);
  total_sum <= total_sum + cache[3039];
endrule
rule s3041(sum_count == 3041);
  total_sum <= total_sum + cache[3040];
endrule
rule s3042(sum_count == 3042);
  total_sum <= total_sum + cache[3041];
endrule
rule s3043(sum_count == 3043);
  total_sum <= total_sum + cache[3042];
endrule
rule s3044(sum_count == 3044);
  total_sum <= total_sum + cache[3043];
endrule
rule s3045(sum_count == 3045);
  total_sum <= total_sum + cache[3044];
endrule
rule s3046(sum_count == 3046);
  total_sum <= total_sum + cache[3045];
endrule
rule s3047(sum_count == 3047);
  total_sum <= total_sum + cache[3046];
endrule
rule s3048(sum_count == 3048);
  total_sum <= total_sum + cache[3047];
endrule
rule s3049(sum_count == 3049);
  total_sum <= total_sum + cache[3048];
endrule
rule s3050(sum_count == 3050);
  total_sum <= total_sum + cache[3049];
endrule
rule s3051(sum_count == 3051);
  total_sum <= total_sum + cache[3050];
endrule
rule s3052(sum_count == 3052);
  total_sum <= total_sum + cache[3051];
endrule
rule s3053(sum_count == 3053);
  total_sum <= total_sum + cache[3052];
endrule
rule s3054(sum_count == 3054);
  total_sum <= total_sum + cache[3053];
endrule
rule s3055(sum_count == 3055);
  total_sum <= total_sum + cache[3054];
endrule
rule s3056(sum_count == 3056);
  total_sum <= total_sum + cache[3055];
endrule
rule s3057(sum_count == 3057);
  total_sum <= total_sum + cache[3056];
endrule
rule s3058(sum_count == 3058);
  total_sum <= total_sum + cache[3057];
endrule
rule s3059(sum_count == 3059);
  total_sum <= total_sum + cache[3058];
endrule
rule s3060(sum_count == 3060);
  total_sum <= total_sum + cache[3059];
endrule
rule s3061(sum_count == 3061);
  total_sum <= total_sum + cache[3060];
endrule
rule s3062(sum_count == 3062);
  total_sum <= total_sum + cache[3061];
endrule
rule s3063(sum_count == 3063);
  total_sum <= total_sum + cache[3062];
endrule
rule s3064(sum_count == 3064);
  total_sum <= total_sum + cache[3063];
endrule
rule s3065(sum_count == 3065);
  total_sum <= total_sum + cache[3064];
endrule
rule s3066(sum_count == 3066);
  total_sum <= total_sum + cache[3065];
endrule
rule s3067(sum_count == 3067);
  total_sum <= total_sum + cache[3066];
endrule
rule s3068(sum_count == 3068);
  total_sum <= total_sum + cache[3067];
endrule
rule s3069(sum_count == 3069);
  total_sum <= total_sum + cache[3068];
endrule
rule s3070(sum_count == 3070);
  total_sum <= total_sum + cache[3069];
endrule
rule s3071(sum_count == 3071);
  total_sum <= total_sum + cache[3070];
endrule
rule s3072(sum_count == 3072);
  total_sum <= total_sum + cache[3071];
endrule
rule s3073(sum_count == 3073);
  total_sum <= total_sum + cache[3072];
endrule
rule s3074(sum_count == 3074);
  total_sum <= total_sum + cache[3073];
endrule
rule s3075(sum_count == 3075);
  total_sum <= total_sum + cache[3074];
endrule
rule s3076(sum_count == 3076);
  total_sum <= total_sum + cache[3075];
endrule
rule s3077(sum_count == 3077);
  total_sum <= total_sum + cache[3076];
endrule
rule s3078(sum_count == 3078);
  total_sum <= total_sum + cache[3077];
endrule
rule s3079(sum_count == 3079);
  total_sum <= total_sum + cache[3078];
endrule
rule s3080(sum_count == 3080);
  total_sum <= total_sum + cache[3079];
endrule
rule s3081(sum_count == 3081);
  total_sum <= total_sum + cache[3080];
endrule
rule s3082(sum_count == 3082);
  total_sum <= total_sum + cache[3081];
endrule
rule s3083(sum_count == 3083);
  total_sum <= total_sum + cache[3082];
endrule
rule s3084(sum_count == 3084);
  total_sum <= total_sum + cache[3083];
endrule
rule s3085(sum_count == 3085);
  total_sum <= total_sum + cache[3084];
endrule
rule s3086(sum_count == 3086);
  total_sum <= total_sum + cache[3085];
endrule
rule s3087(sum_count == 3087);
  total_sum <= total_sum + cache[3086];
endrule
rule s3088(sum_count == 3088);
  total_sum <= total_sum + cache[3087];
endrule
rule s3089(sum_count == 3089);
  total_sum <= total_sum + cache[3088];
endrule
rule s3090(sum_count == 3090);
  total_sum <= total_sum + cache[3089];
endrule
rule s3091(sum_count == 3091);
  total_sum <= total_sum + cache[3090];
endrule
rule s3092(sum_count == 3092);
  total_sum <= total_sum + cache[3091];
endrule
rule s3093(sum_count == 3093);
  total_sum <= total_sum + cache[3092];
endrule
rule s3094(sum_count == 3094);
  total_sum <= total_sum + cache[3093];
endrule
rule s3095(sum_count == 3095);
  total_sum <= total_sum + cache[3094];
endrule
rule s3096(sum_count == 3096);
  total_sum <= total_sum + cache[3095];
endrule
rule s3097(sum_count == 3097);
  total_sum <= total_sum + cache[3096];
endrule
rule s3098(sum_count == 3098);
  total_sum <= total_sum + cache[3097];
endrule
rule s3099(sum_count == 3099);
  total_sum <= total_sum + cache[3098];
endrule
rule s3100(sum_count == 3100);
  total_sum <= total_sum + cache[3099];
endrule
rule s3101(sum_count == 3101);
  total_sum <= total_sum + cache[3100];
endrule
rule s3102(sum_count == 3102);
  total_sum <= total_sum + cache[3101];
endrule
rule s3103(sum_count == 3103);
  total_sum <= total_sum + cache[3102];
endrule
rule s3104(sum_count == 3104);
  total_sum <= total_sum + cache[3103];
endrule
rule s3105(sum_count == 3105);
  total_sum <= total_sum + cache[3104];
endrule
rule s3106(sum_count == 3106);
  total_sum <= total_sum + cache[3105];
endrule
rule s3107(sum_count == 3107);
  total_sum <= total_sum + cache[3106];
endrule
rule s3108(sum_count == 3108);
  total_sum <= total_sum + cache[3107];
endrule
rule s3109(sum_count == 3109);
  total_sum <= total_sum + cache[3108];
endrule
rule s3110(sum_count == 3110);
  total_sum <= total_sum + cache[3109];
endrule
rule s3111(sum_count == 3111);
  total_sum <= total_sum + cache[3110];
endrule
rule s3112(sum_count == 3112);
  total_sum <= total_sum + cache[3111];
endrule
rule s3113(sum_count == 3113);
  total_sum <= total_sum + cache[3112];
endrule
rule s3114(sum_count == 3114);
  total_sum <= total_sum + cache[3113];
endrule
rule s3115(sum_count == 3115);
  total_sum <= total_sum + cache[3114];
endrule
rule s3116(sum_count == 3116);
  total_sum <= total_sum + cache[3115];
endrule
rule s3117(sum_count == 3117);
  total_sum <= total_sum + cache[3116];
endrule
rule s3118(sum_count == 3118);
  total_sum <= total_sum + cache[3117];
endrule
rule s3119(sum_count == 3119);
  total_sum <= total_sum + cache[3118];
endrule
rule s3120(sum_count == 3120);
  total_sum <= total_sum + cache[3119];
endrule
rule s3121(sum_count == 3121);
  total_sum <= total_sum + cache[3120];
endrule
rule s3122(sum_count == 3122);
  total_sum <= total_sum + cache[3121];
endrule
rule s3123(sum_count == 3123);
  total_sum <= total_sum + cache[3122];
endrule
rule s3124(sum_count == 3124);
  total_sum <= total_sum + cache[3123];
endrule
rule s3125(sum_count == 3125);
  total_sum <= total_sum + cache[3124];
endrule
rule s3126(sum_count == 3126);
  total_sum <= total_sum + cache[3125];
endrule
rule s3127(sum_count == 3127);
  total_sum <= total_sum + cache[3126];
endrule
rule s3128(sum_count == 3128);
  total_sum <= total_sum + cache[3127];
endrule
rule s3129(sum_count == 3129);
  total_sum <= total_sum + cache[3128];
endrule
rule s3130(sum_count == 3130);
  total_sum <= total_sum + cache[3129];
endrule
rule s3131(sum_count == 3131);
  total_sum <= total_sum + cache[3130];
endrule
rule s3132(sum_count == 3132);
  total_sum <= total_sum + cache[3131];
endrule
rule s3133(sum_count == 3133);
  total_sum <= total_sum + cache[3132];
endrule
rule s3134(sum_count == 3134);
  total_sum <= total_sum + cache[3133];
endrule
rule s3135(sum_count == 3135);
  total_sum <= total_sum + cache[3134];
endrule
rule s3136(sum_count == 3136);
  total_sum <= total_sum + cache[3135];
endrule
rule s3137(sum_count == 3137);
  total_sum <= total_sum + cache[3136];
endrule
rule s3138(sum_count == 3138);
  total_sum <= total_sum + cache[3137];
endrule
rule s3139(sum_count == 3139);
  total_sum <= total_sum + cache[3138];
endrule
rule s3140(sum_count == 3140);
  total_sum <= total_sum + cache[3139];
endrule
rule s3141(sum_count == 3141);
  total_sum <= total_sum + cache[3140];
endrule
rule s3142(sum_count == 3142);
  total_sum <= total_sum + cache[3141];
endrule
rule s3143(sum_count == 3143);
  total_sum <= total_sum + cache[3142];
endrule
rule s3144(sum_count == 3144);
  total_sum <= total_sum + cache[3143];
endrule
rule s3145(sum_count == 3145);
  total_sum <= total_sum + cache[3144];
endrule
rule s3146(sum_count == 3146);
  total_sum <= total_sum + cache[3145];
endrule
rule s3147(sum_count == 3147);
  total_sum <= total_sum + cache[3146];
endrule
rule s3148(sum_count == 3148);
  total_sum <= total_sum + cache[3147];
endrule
rule s3149(sum_count == 3149);
  total_sum <= total_sum + cache[3148];
endrule
rule s3150(sum_count == 3150);
  total_sum <= total_sum + cache[3149];
endrule
rule s3151(sum_count == 3151);
  total_sum <= total_sum + cache[3150];
endrule
rule s3152(sum_count == 3152);
  total_sum <= total_sum + cache[3151];
endrule
rule s3153(sum_count == 3153);
  total_sum <= total_sum + cache[3152];
endrule
rule s3154(sum_count == 3154);
  total_sum <= total_sum + cache[3153];
endrule
rule s3155(sum_count == 3155);
  total_sum <= total_sum + cache[3154];
endrule
rule s3156(sum_count == 3156);
  total_sum <= total_sum + cache[3155];
endrule
rule s3157(sum_count == 3157);
  total_sum <= total_sum + cache[3156];
endrule
rule s3158(sum_count == 3158);
  total_sum <= total_sum + cache[3157];
endrule
rule s3159(sum_count == 3159);
  total_sum <= total_sum + cache[3158];
endrule
rule s3160(sum_count == 3160);
  total_sum <= total_sum + cache[3159];
endrule
rule s3161(sum_count == 3161);
  total_sum <= total_sum + cache[3160];
endrule
rule s3162(sum_count == 3162);
  total_sum <= total_sum + cache[3161];
endrule
rule s3163(sum_count == 3163);
  total_sum <= total_sum + cache[3162];
endrule
rule s3164(sum_count == 3164);
  total_sum <= total_sum + cache[3163];
endrule
rule s3165(sum_count == 3165);
  total_sum <= total_sum + cache[3164];
endrule
rule s3166(sum_count == 3166);
  total_sum <= total_sum + cache[3165];
endrule
rule s3167(sum_count == 3167);
  total_sum <= total_sum + cache[3166];
endrule
rule s3168(sum_count == 3168);
  total_sum <= total_sum + cache[3167];
endrule
rule s3169(sum_count == 3169);
  total_sum <= total_sum + cache[3168];
endrule
rule s3170(sum_count == 3170);
  total_sum <= total_sum + cache[3169];
endrule
rule s3171(sum_count == 3171);
  total_sum <= total_sum + cache[3170];
endrule
rule s3172(sum_count == 3172);
  total_sum <= total_sum + cache[3171];
endrule
rule s3173(sum_count == 3173);
  total_sum <= total_sum + cache[3172];
endrule
rule s3174(sum_count == 3174);
  total_sum <= total_sum + cache[3173];
endrule
rule s3175(sum_count == 3175);
  total_sum <= total_sum + cache[3174];
endrule
rule s3176(sum_count == 3176);
  total_sum <= total_sum + cache[3175];
endrule
rule s3177(sum_count == 3177);
  total_sum <= total_sum + cache[3176];
endrule
rule s3178(sum_count == 3178);
  total_sum <= total_sum + cache[3177];
endrule
rule s3179(sum_count == 3179);
  total_sum <= total_sum + cache[3178];
endrule
rule s3180(sum_count == 3180);
  total_sum <= total_sum + cache[3179];
endrule
rule s3181(sum_count == 3181);
  total_sum <= total_sum + cache[3180];
endrule
rule s3182(sum_count == 3182);
  total_sum <= total_sum + cache[3181];
endrule
rule s3183(sum_count == 3183);
  total_sum <= total_sum + cache[3182];
endrule
rule s3184(sum_count == 3184);
  total_sum <= total_sum + cache[3183];
endrule
rule s3185(sum_count == 3185);
  total_sum <= total_sum + cache[3184];
endrule
rule s3186(sum_count == 3186);
  total_sum <= total_sum + cache[3185];
endrule
rule s3187(sum_count == 3187);
  total_sum <= total_sum + cache[3186];
endrule
rule s3188(sum_count == 3188);
  total_sum <= total_sum + cache[3187];
endrule
rule s3189(sum_count == 3189);
  total_sum <= total_sum + cache[3188];
endrule
rule s3190(sum_count == 3190);
  total_sum <= total_sum + cache[3189];
endrule
rule s3191(sum_count == 3191);
  total_sum <= total_sum + cache[3190];
endrule
rule s3192(sum_count == 3192);
  total_sum <= total_sum + cache[3191];
endrule
rule s3193(sum_count == 3193);
  total_sum <= total_sum + cache[3192];
endrule
rule s3194(sum_count == 3194);
  total_sum <= total_sum + cache[3193];
endrule
rule s3195(sum_count == 3195);
  total_sum <= total_sum + cache[3194];
endrule
rule s3196(sum_count == 3196);
  total_sum <= total_sum + cache[3195];
endrule
rule s3197(sum_count == 3197);
  total_sum <= total_sum + cache[3196];
endrule
rule s3198(sum_count == 3198);
  total_sum <= total_sum + cache[3197];
endrule
rule s3199(sum_count == 3199);
  total_sum <= total_sum + cache[3198];
endrule
rule s3200(sum_count == 3200);
  total_sum <= total_sum + cache[3199];
endrule
rule s3201(sum_count == 3201);
  total_sum <= total_sum + cache[3200];
endrule
rule s3202(sum_count == 3202);
  total_sum <= total_sum + cache[3201];
endrule
rule s3203(sum_count == 3203);
  total_sum <= total_sum + cache[3202];
endrule
rule s3204(sum_count == 3204);
  total_sum <= total_sum + cache[3203];
endrule
rule s3205(sum_count == 3205);
  total_sum <= total_sum + cache[3204];
endrule
rule s3206(sum_count == 3206);
  total_sum <= total_sum + cache[3205];
endrule
rule s3207(sum_count == 3207);
  total_sum <= total_sum + cache[3206];
endrule
rule s3208(sum_count == 3208);
  total_sum <= total_sum + cache[3207];
endrule
rule s3209(sum_count == 3209);
  total_sum <= total_sum + cache[3208];
endrule
rule s3210(sum_count == 3210);
  total_sum <= total_sum + cache[3209];
endrule
rule s3211(sum_count == 3211);
  total_sum <= total_sum + cache[3210];
endrule
rule s3212(sum_count == 3212);
  total_sum <= total_sum + cache[3211];
endrule
rule s3213(sum_count == 3213);
  total_sum <= total_sum + cache[3212];
endrule
rule s3214(sum_count == 3214);
  total_sum <= total_sum + cache[3213];
endrule
rule s3215(sum_count == 3215);
  total_sum <= total_sum + cache[3214];
endrule
rule s3216(sum_count == 3216);
  total_sum <= total_sum + cache[3215];
endrule
rule s3217(sum_count == 3217);
  total_sum <= total_sum + cache[3216];
endrule
rule s3218(sum_count == 3218);
  total_sum <= total_sum + cache[3217];
endrule
rule s3219(sum_count == 3219);
  total_sum <= total_sum + cache[3218];
endrule
rule s3220(sum_count == 3220);
  total_sum <= total_sum + cache[3219];
endrule
rule s3221(sum_count == 3221);
  total_sum <= total_sum + cache[3220];
endrule
rule s3222(sum_count == 3222);
  total_sum <= total_sum + cache[3221];
endrule
rule s3223(sum_count == 3223);
  total_sum <= total_sum + cache[3222];
endrule
rule s3224(sum_count == 3224);
  total_sum <= total_sum + cache[3223];
endrule
rule s3225(sum_count == 3225);
  total_sum <= total_sum + cache[3224];
endrule
rule s3226(sum_count == 3226);
  total_sum <= total_sum + cache[3225];
endrule
rule s3227(sum_count == 3227);
  total_sum <= total_sum + cache[3226];
endrule
rule s3228(sum_count == 3228);
  total_sum <= total_sum + cache[3227];
endrule
rule s3229(sum_count == 3229);
  total_sum <= total_sum + cache[3228];
endrule
rule s3230(sum_count == 3230);
  total_sum <= total_sum + cache[3229];
endrule
rule s3231(sum_count == 3231);
  total_sum <= total_sum + cache[3230];
endrule
rule s3232(sum_count == 3232);
  total_sum <= total_sum + cache[3231];
endrule
rule s3233(sum_count == 3233);
  total_sum <= total_sum + cache[3232];
endrule
rule s3234(sum_count == 3234);
  total_sum <= total_sum + cache[3233];
endrule
rule s3235(sum_count == 3235);
  total_sum <= total_sum + cache[3234];
endrule
rule s3236(sum_count == 3236);
  total_sum <= total_sum + cache[3235];
endrule
rule s3237(sum_count == 3237);
  total_sum <= total_sum + cache[3236];
endrule
rule s3238(sum_count == 3238);
  total_sum <= total_sum + cache[3237];
endrule
rule s3239(sum_count == 3239);
  total_sum <= total_sum + cache[3238];
endrule
rule s3240(sum_count == 3240);
  total_sum <= total_sum + cache[3239];
endrule
rule s3241(sum_count == 3241);
  total_sum <= total_sum + cache[3240];
endrule
rule s3242(sum_count == 3242);
  total_sum <= total_sum + cache[3241];
endrule
rule s3243(sum_count == 3243);
  total_sum <= total_sum + cache[3242];
endrule
rule s3244(sum_count == 3244);
  total_sum <= total_sum + cache[3243];
endrule
rule s3245(sum_count == 3245);
  total_sum <= total_sum + cache[3244];
endrule
rule s3246(sum_count == 3246);
  total_sum <= total_sum + cache[3245];
endrule
rule s3247(sum_count == 3247);
  total_sum <= total_sum + cache[3246];
endrule
rule s3248(sum_count == 3248);
  total_sum <= total_sum + cache[3247];
endrule
rule s3249(sum_count == 3249);
  total_sum <= total_sum + cache[3248];
endrule
rule s3250(sum_count == 3250);
  total_sum <= total_sum + cache[3249];
endrule
rule s3251(sum_count == 3251);
  total_sum <= total_sum + cache[3250];
endrule
rule s3252(sum_count == 3252);
  total_sum <= total_sum + cache[3251];
endrule
rule s3253(sum_count == 3253);
  total_sum <= total_sum + cache[3252];
endrule
rule s3254(sum_count == 3254);
  total_sum <= total_sum + cache[3253];
endrule
rule s3255(sum_count == 3255);
  total_sum <= total_sum + cache[3254];
endrule
rule s3256(sum_count == 3256);
  total_sum <= total_sum + cache[3255];
endrule
rule s3257(sum_count == 3257);
  total_sum <= total_sum + cache[3256];
endrule
rule s3258(sum_count == 3258);
  total_sum <= total_sum + cache[3257];
endrule
rule s3259(sum_count == 3259);
  total_sum <= total_sum + cache[3258];
endrule
rule s3260(sum_count == 3260);
  total_sum <= total_sum + cache[3259];
endrule
rule s3261(sum_count == 3261);
  total_sum <= total_sum + cache[3260];
endrule
rule s3262(sum_count == 3262);
  total_sum <= total_sum + cache[3261];
endrule
rule s3263(sum_count == 3263);
  total_sum <= total_sum + cache[3262];
endrule
rule s3264(sum_count == 3264);
  total_sum <= total_sum + cache[3263];
endrule
rule s3265(sum_count == 3265);
  total_sum <= total_sum + cache[3264];
endrule
rule s3266(sum_count == 3266);
  total_sum <= total_sum + cache[3265];
endrule
rule s3267(sum_count == 3267);
  total_sum <= total_sum + cache[3266];
endrule
rule s3268(sum_count == 3268);
  total_sum <= total_sum + cache[3267];
endrule
rule s3269(sum_count == 3269);
  total_sum <= total_sum + cache[3268];
endrule
rule s3270(sum_count == 3270);
  total_sum <= total_sum + cache[3269];
endrule
rule s3271(sum_count == 3271);
  total_sum <= total_sum + cache[3270];
endrule
rule s3272(sum_count == 3272);
  total_sum <= total_sum + cache[3271];
endrule
rule s3273(sum_count == 3273);
  total_sum <= total_sum + cache[3272];
endrule
rule s3274(sum_count == 3274);
  total_sum <= total_sum + cache[3273];
endrule
rule s3275(sum_count == 3275);
  total_sum <= total_sum + cache[3274];
endrule
rule s3276(sum_count == 3276);
  total_sum <= total_sum + cache[3275];
endrule
rule s3277(sum_count == 3277);
  total_sum <= total_sum + cache[3276];
endrule
rule s3278(sum_count == 3278);
  total_sum <= total_sum + cache[3277];
endrule
rule s3279(sum_count == 3279);
  total_sum <= total_sum + cache[3278];
endrule
rule s3280(sum_count == 3280);
  total_sum <= total_sum + cache[3279];
endrule
rule s3281(sum_count == 3281);
  total_sum <= total_sum + cache[3280];
endrule
rule s3282(sum_count == 3282);
  total_sum <= total_sum + cache[3281];
endrule
rule s3283(sum_count == 3283);
  total_sum <= total_sum + cache[3282];
endrule
rule s3284(sum_count == 3284);
  total_sum <= total_sum + cache[3283];
endrule
rule s3285(sum_count == 3285);
  total_sum <= total_sum + cache[3284];
endrule
rule s3286(sum_count == 3286);
  total_sum <= total_sum + cache[3285];
endrule
rule s3287(sum_count == 3287);
  total_sum <= total_sum + cache[3286];
endrule
rule s3288(sum_count == 3288);
  total_sum <= total_sum + cache[3287];
endrule
rule s3289(sum_count == 3289);
  total_sum <= total_sum + cache[3288];
endrule
rule s3290(sum_count == 3290);
  total_sum <= total_sum + cache[3289];
endrule
rule s3291(sum_count == 3291);
  total_sum <= total_sum + cache[3290];
endrule
rule s3292(sum_count == 3292);
  total_sum <= total_sum + cache[3291];
endrule
rule s3293(sum_count == 3293);
  total_sum <= total_sum + cache[3292];
endrule
rule s3294(sum_count == 3294);
  total_sum <= total_sum + cache[3293];
endrule
rule s3295(sum_count == 3295);
  total_sum <= total_sum + cache[3294];
endrule
rule s3296(sum_count == 3296);
  total_sum <= total_sum + cache[3295];
endrule
rule s3297(sum_count == 3297);
  total_sum <= total_sum + cache[3296];
endrule
rule s3298(sum_count == 3298);
  total_sum <= total_sum + cache[3297];
endrule
rule s3299(sum_count == 3299);
  total_sum <= total_sum + cache[3298];
endrule
rule s3300(sum_count == 3300);
  total_sum <= total_sum + cache[3299];
endrule
rule s3301(sum_count == 3301);
  total_sum <= total_sum + cache[3300];
endrule
rule s3302(sum_count == 3302);
  total_sum <= total_sum + cache[3301];
endrule
rule s3303(sum_count == 3303);
  total_sum <= total_sum + cache[3302];
endrule
rule s3304(sum_count == 3304);
  total_sum <= total_sum + cache[3303];
endrule
rule s3305(sum_count == 3305);
  total_sum <= total_sum + cache[3304];
endrule
rule s3306(sum_count == 3306);
  total_sum <= total_sum + cache[3305];
endrule
rule s3307(sum_count == 3307);
  total_sum <= total_sum + cache[3306];
endrule
rule s3308(sum_count == 3308);
  total_sum <= total_sum + cache[3307];
endrule
rule s3309(sum_count == 3309);
  total_sum <= total_sum + cache[3308];
endrule
rule s3310(sum_count == 3310);
  total_sum <= total_sum + cache[3309];
endrule
rule s3311(sum_count == 3311);
  total_sum <= total_sum + cache[3310];
endrule
rule s3312(sum_count == 3312);
  total_sum <= total_sum + cache[3311];
endrule
rule s3313(sum_count == 3313);
  total_sum <= total_sum + cache[3312];
endrule
rule s3314(sum_count == 3314);
  total_sum <= total_sum + cache[3313];
endrule
rule s3315(sum_count == 3315);
  total_sum <= total_sum + cache[3314];
endrule
rule s3316(sum_count == 3316);
  total_sum <= total_sum + cache[3315];
endrule
rule s3317(sum_count == 3317);
  total_sum <= total_sum + cache[3316];
endrule
rule s3318(sum_count == 3318);
  total_sum <= total_sum + cache[3317];
endrule
rule s3319(sum_count == 3319);
  total_sum <= total_sum + cache[3318];
endrule
rule s3320(sum_count == 3320);
  total_sum <= total_sum + cache[3319];
endrule
rule s3321(sum_count == 3321);
  total_sum <= total_sum + cache[3320];
endrule
rule s3322(sum_count == 3322);
  total_sum <= total_sum + cache[3321];
endrule
rule s3323(sum_count == 3323);
  total_sum <= total_sum + cache[3322];
endrule
rule s3324(sum_count == 3324);
  total_sum <= total_sum + cache[3323];
endrule
rule s3325(sum_count == 3325);
  total_sum <= total_sum + cache[3324];
endrule
rule s3326(sum_count == 3326);
  total_sum <= total_sum + cache[3325];
endrule
rule s3327(sum_count == 3327);
  total_sum <= total_sum + cache[3326];
endrule
rule s3328(sum_count == 3328);
  total_sum <= total_sum + cache[3327];
endrule
rule s3329(sum_count == 3329);
  total_sum <= total_sum + cache[3328];
endrule
rule s3330(sum_count == 3330);
  total_sum <= total_sum + cache[3329];
endrule
rule s3331(sum_count == 3331);
  total_sum <= total_sum + cache[3330];
endrule
rule s3332(sum_count == 3332);
  total_sum <= total_sum + cache[3331];
endrule
rule s3333(sum_count == 3333);
  total_sum <= total_sum + cache[3332];
endrule
rule s3334(sum_count == 3334);
  total_sum <= total_sum + cache[3333];
endrule
rule s3335(sum_count == 3335);
  total_sum <= total_sum + cache[3334];
endrule
rule s3336(sum_count == 3336);
  total_sum <= total_sum + cache[3335];
endrule
rule s3337(sum_count == 3337);
  total_sum <= total_sum + cache[3336];
endrule
rule s3338(sum_count == 3338);
  total_sum <= total_sum + cache[3337];
endrule
rule s3339(sum_count == 3339);
  total_sum <= total_sum + cache[3338];
endrule
rule s3340(sum_count == 3340);
  total_sum <= total_sum + cache[3339];
endrule
rule s3341(sum_count == 3341);
  total_sum <= total_sum + cache[3340];
endrule
rule s3342(sum_count == 3342);
  total_sum <= total_sum + cache[3341];
endrule
rule s3343(sum_count == 3343);
  total_sum <= total_sum + cache[3342];
endrule
rule s3344(sum_count == 3344);
  total_sum <= total_sum + cache[3343];
endrule
rule s3345(sum_count == 3345);
  total_sum <= total_sum + cache[3344];
endrule
rule s3346(sum_count == 3346);
  total_sum <= total_sum + cache[3345];
endrule
rule s3347(sum_count == 3347);
  total_sum <= total_sum + cache[3346];
endrule
rule s3348(sum_count == 3348);
  total_sum <= total_sum + cache[3347];
endrule
rule s3349(sum_count == 3349);
  total_sum <= total_sum + cache[3348];
endrule
rule s3350(sum_count == 3350);
  total_sum <= total_sum + cache[3349];
endrule
rule s3351(sum_count == 3351);
  total_sum <= total_sum + cache[3350];
endrule
rule s3352(sum_count == 3352);
  total_sum <= total_sum + cache[3351];
endrule
rule s3353(sum_count == 3353);
  total_sum <= total_sum + cache[3352];
endrule
rule s3354(sum_count == 3354);
  total_sum <= total_sum + cache[3353];
endrule
rule s3355(sum_count == 3355);
  total_sum <= total_sum + cache[3354];
endrule
rule s3356(sum_count == 3356);
  total_sum <= total_sum + cache[3355];
endrule
rule s3357(sum_count == 3357);
  total_sum <= total_sum + cache[3356];
endrule
rule s3358(sum_count == 3358);
  total_sum <= total_sum + cache[3357];
endrule
rule s3359(sum_count == 3359);
  total_sum <= total_sum + cache[3358];
endrule
rule s3360(sum_count == 3360);
  total_sum <= total_sum + cache[3359];
endrule
rule s3361(sum_count == 3361);
  total_sum <= total_sum + cache[3360];
endrule
rule s3362(sum_count == 3362);
  total_sum <= total_sum + cache[3361];
endrule
rule s3363(sum_count == 3363);
  total_sum <= total_sum + cache[3362];
endrule
rule s3364(sum_count == 3364);
  total_sum <= total_sum + cache[3363];
endrule
rule s3365(sum_count == 3365);
  total_sum <= total_sum + cache[3364];
endrule
rule s3366(sum_count == 3366);
  total_sum <= total_sum + cache[3365];
endrule
rule s3367(sum_count == 3367);
  total_sum <= total_sum + cache[3366];
endrule
rule s3368(sum_count == 3368);
  total_sum <= total_sum + cache[3367];
endrule
rule s3369(sum_count == 3369);
  total_sum <= total_sum + cache[3368];
endrule
rule s3370(sum_count == 3370);
  total_sum <= total_sum + cache[3369];
endrule
rule s3371(sum_count == 3371);
  total_sum <= total_sum + cache[3370];
endrule
rule s3372(sum_count == 3372);
  total_sum <= total_sum + cache[3371];
endrule
rule s3373(sum_count == 3373);
  total_sum <= total_sum + cache[3372];
endrule
rule s3374(sum_count == 3374);
  total_sum <= total_sum + cache[3373];
endrule
rule s3375(sum_count == 3375);
  total_sum <= total_sum + cache[3374];
endrule
rule s3376(sum_count == 3376);
  total_sum <= total_sum + cache[3375];
endrule
rule s3377(sum_count == 3377);
  total_sum <= total_sum + cache[3376];
endrule
rule s3378(sum_count == 3378);
  total_sum <= total_sum + cache[3377];
endrule
rule s3379(sum_count == 3379);
  total_sum <= total_sum + cache[3378];
endrule
rule s3380(sum_count == 3380);
  total_sum <= total_sum + cache[3379];
endrule
rule s3381(sum_count == 3381);
  total_sum <= total_sum + cache[3380];
endrule
rule s3382(sum_count == 3382);
  total_sum <= total_sum + cache[3381];
endrule
rule s3383(sum_count == 3383);
  total_sum <= total_sum + cache[3382];
endrule
rule s3384(sum_count == 3384);
  total_sum <= total_sum + cache[3383];
endrule
rule s3385(sum_count == 3385);
  total_sum <= total_sum + cache[3384];
endrule
rule s3386(sum_count == 3386);
  total_sum <= total_sum + cache[3385];
endrule
rule s3387(sum_count == 3387);
  total_sum <= total_sum + cache[3386];
endrule
rule s3388(sum_count == 3388);
  total_sum <= total_sum + cache[3387];
endrule
rule s3389(sum_count == 3389);
  total_sum <= total_sum + cache[3388];
endrule
rule s3390(sum_count == 3390);
  total_sum <= total_sum + cache[3389];
endrule
rule s3391(sum_count == 3391);
  total_sum <= total_sum + cache[3390];
endrule
rule s3392(sum_count == 3392);
  total_sum <= total_sum + cache[3391];
endrule
rule s3393(sum_count == 3393);
  total_sum <= total_sum + cache[3392];
endrule
rule s3394(sum_count == 3394);
  total_sum <= total_sum + cache[3393];
endrule
rule s3395(sum_count == 3395);
  total_sum <= total_sum + cache[3394];
endrule
rule s3396(sum_count == 3396);
  total_sum <= total_sum + cache[3395];
endrule
rule s3397(sum_count == 3397);
  total_sum <= total_sum + cache[3396];
endrule
rule s3398(sum_count == 3398);
  total_sum <= total_sum + cache[3397];
endrule
rule s3399(sum_count == 3399);
  total_sum <= total_sum + cache[3398];
endrule
rule s3400(sum_count == 3400);
  total_sum <= total_sum + cache[3399];
endrule
rule s3401(sum_count == 3401);
  total_sum <= total_sum + cache[3400];
endrule
rule s3402(sum_count == 3402);
  total_sum <= total_sum + cache[3401];
endrule
rule s3403(sum_count == 3403);
  total_sum <= total_sum + cache[3402];
endrule
rule s3404(sum_count == 3404);
  total_sum <= total_sum + cache[3403];
endrule
rule s3405(sum_count == 3405);
  total_sum <= total_sum + cache[3404];
endrule
rule s3406(sum_count == 3406);
  total_sum <= total_sum + cache[3405];
endrule
rule s3407(sum_count == 3407);
  total_sum <= total_sum + cache[3406];
endrule
rule s3408(sum_count == 3408);
  total_sum <= total_sum + cache[3407];
endrule
rule s3409(sum_count == 3409);
  total_sum <= total_sum + cache[3408];
endrule
rule s3410(sum_count == 3410);
  total_sum <= total_sum + cache[3409];
endrule
rule s3411(sum_count == 3411);
  total_sum <= total_sum + cache[3410];
endrule
rule s3412(sum_count == 3412);
  total_sum <= total_sum + cache[3411];
endrule
rule s3413(sum_count == 3413);
  total_sum <= total_sum + cache[3412];
endrule
rule s3414(sum_count == 3414);
  total_sum <= total_sum + cache[3413];
endrule
rule s3415(sum_count == 3415);
  total_sum <= total_sum + cache[3414];
endrule
rule s3416(sum_count == 3416);
  total_sum <= total_sum + cache[3415];
endrule
rule s3417(sum_count == 3417);
  total_sum <= total_sum + cache[3416];
endrule
rule s3418(sum_count == 3418);
  total_sum <= total_sum + cache[3417];
endrule
rule s3419(sum_count == 3419);
  total_sum <= total_sum + cache[3418];
endrule
rule s3420(sum_count == 3420);
  total_sum <= total_sum + cache[3419];
endrule
rule s3421(sum_count == 3421);
  total_sum <= total_sum + cache[3420];
endrule
rule s3422(sum_count == 3422);
  total_sum <= total_sum + cache[3421];
endrule
rule s3423(sum_count == 3423);
  total_sum <= total_sum + cache[3422];
endrule
rule s3424(sum_count == 3424);
  total_sum <= total_sum + cache[3423];
endrule
rule s3425(sum_count == 3425);
  total_sum <= total_sum + cache[3424];
endrule
rule s3426(sum_count == 3426);
  total_sum <= total_sum + cache[3425];
endrule
rule s3427(sum_count == 3427);
  total_sum <= total_sum + cache[3426];
endrule
rule s3428(sum_count == 3428);
  total_sum <= total_sum + cache[3427];
endrule
rule s3429(sum_count == 3429);
  total_sum <= total_sum + cache[3428];
endrule
rule s3430(sum_count == 3430);
  total_sum <= total_sum + cache[3429];
endrule
rule s3431(sum_count == 3431);
  total_sum <= total_sum + cache[3430];
endrule
rule s3432(sum_count == 3432);
  total_sum <= total_sum + cache[3431];
endrule
rule s3433(sum_count == 3433);
  total_sum <= total_sum + cache[3432];
endrule
rule s3434(sum_count == 3434);
  total_sum <= total_sum + cache[3433];
endrule
rule s3435(sum_count == 3435);
  total_sum <= total_sum + cache[3434];
endrule
rule s3436(sum_count == 3436);
  total_sum <= total_sum + cache[3435];
endrule
rule s3437(sum_count == 3437);
  total_sum <= total_sum + cache[3436];
endrule
rule s3438(sum_count == 3438);
  total_sum <= total_sum + cache[3437];
endrule
rule s3439(sum_count == 3439);
  total_sum <= total_sum + cache[3438];
endrule
rule s3440(sum_count == 3440);
  total_sum <= total_sum + cache[3439];
endrule
rule s3441(sum_count == 3441);
  total_sum <= total_sum + cache[3440];
endrule
rule s3442(sum_count == 3442);
  total_sum <= total_sum + cache[3441];
endrule
rule s3443(sum_count == 3443);
  total_sum <= total_sum + cache[3442];
endrule
rule s3444(sum_count == 3444);
  total_sum <= total_sum + cache[3443];
endrule
rule s3445(sum_count == 3445);
  total_sum <= total_sum + cache[3444];
endrule
rule s3446(sum_count == 3446);
  total_sum <= total_sum + cache[3445];
endrule
rule s3447(sum_count == 3447);
  total_sum <= total_sum + cache[3446];
endrule
rule s3448(sum_count == 3448);
  total_sum <= total_sum + cache[3447];
endrule
rule s3449(sum_count == 3449);
  total_sum <= total_sum + cache[3448];
endrule
rule s3450(sum_count == 3450);
  total_sum <= total_sum + cache[3449];
endrule
rule s3451(sum_count == 3451);
  total_sum <= total_sum + cache[3450];
endrule
rule s3452(sum_count == 3452);
  total_sum <= total_sum + cache[3451];
endrule
rule s3453(sum_count == 3453);
  total_sum <= total_sum + cache[3452];
endrule
rule s3454(sum_count == 3454);
  total_sum <= total_sum + cache[3453];
endrule
rule s3455(sum_count == 3455);
  total_sum <= total_sum + cache[3454];
endrule
rule s3456(sum_count == 3456);
  total_sum <= total_sum + cache[3455];
endrule
rule s3457(sum_count == 3457);
  total_sum <= total_sum + cache[3456];
endrule
rule s3458(sum_count == 3458);
  total_sum <= total_sum + cache[3457];
endrule
rule s3459(sum_count == 3459);
  total_sum <= total_sum + cache[3458];
endrule
rule s3460(sum_count == 3460);
  total_sum <= total_sum + cache[3459];
endrule
rule s3461(sum_count == 3461);
  total_sum <= total_sum + cache[3460];
endrule
rule s3462(sum_count == 3462);
  total_sum <= total_sum + cache[3461];
endrule
rule s3463(sum_count == 3463);
  total_sum <= total_sum + cache[3462];
endrule
rule s3464(sum_count == 3464);
  total_sum <= total_sum + cache[3463];
endrule
rule s3465(sum_count == 3465);
  total_sum <= total_sum + cache[3464];
endrule
rule s3466(sum_count == 3466);
  total_sum <= total_sum + cache[3465];
endrule
rule s3467(sum_count == 3467);
  total_sum <= total_sum + cache[3466];
endrule
rule s3468(sum_count == 3468);
  total_sum <= total_sum + cache[3467];
endrule
rule s3469(sum_count == 3469);
  total_sum <= total_sum + cache[3468];
endrule
rule s3470(sum_count == 3470);
  total_sum <= total_sum + cache[3469];
endrule
rule s3471(sum_count == 3471);
  total_sum <= total_sum + cache[3470];
endrule
rule s3472(sum_count == 3472);
  total_sum <= total_sum + cache[3471];
endrule
rule s3473(sum_count == 3473);
  total_sum <= total_sum + cache[3472];
endrule
rule s3474(sum_count == 3474);
  total_sum <= total_sum + cache[3473];
endrule
rule s3475(sum_count == 3475);
  total_sum <= total_sum + cache[3474];
endrule
rule s3476(sum_count == 3476);
  total_sum <= total_sum + cache[3475];
endrule
rule s3477(sum_count == 3477);
  total_sum <= total_sum + cache[3476];
endrule
rule s3478(sum_count == 3478);
  total_sum <= total_sum + cache[3477];
endrule
rule s3479(sum_count == 3479);
  total_sum <= total_sum + cache[3478];
endrule
rule s3480(sum_count == 3480);
  total_sum <= total_sum + cache[3479];
endrule
rule s3481(sum_count == 3481);
  total_sum <= total_sum + cache[3480];
endrule
rule s3482(sum_count == 3482);
  total_sum <= total_sum + cache[3481];
endrule
rule s3483(sum_count == 3483);
  total_sum <= total_sum + cache[3482];
endrule
rule s3484(sum_count == 3484);
  total_sum <= total_sum + cache[3483];
endrule
rule s3485(sum_count == 3485);
  total_sum <= total_sum + cache[3484];
endrule
rule s3486(sum_count == 3486);
  total_sum <= total_sum + cache[3485];
endrule
rule s3487(sum_count == 3487);
  total_sum <= total_sum + cache[3486];
endrule
rule s3488(sum_count == 3488);
  total_sum <= total_sum + cache[3487];
endrule
rule s3489(sum_count == 3489);
  total_sum <= total_sum + cache[3488];
endrule
rule s3490(sum_count == 3490);
  total_sum <= total_sum + cache[3489];
endrule
rule s3491(sum_count == 3491);
  total_sum <= total_sum + cache[3490];
endrule
rule s3492(sum_count == 3492);
  total_sum <= total_sum + cache[3491];
endrule
rule s3493(sum_count == 3493);
  total_sum <= total_sum + cache[3492];
endrule
rule s3494(sum_count == 3494);
  total_sum <= total_sum + cache[3493];
endrule
rule s3495(sum_count == 3495);
  total_sum <= total_sum + cache[3494];
endrule
rule s3496(sum_count == 3496);
  total_sum <= total_sum + cache[3495];
endrule
rule s3497(sum_count == 3497);
  total_sum <= total_sum + cache[3496];
endrule
rule s3498(sum_count == 3498);
  total_sum <= total_sum + cache[3497];
endrule
rule s3499(sum_count == 3499);
  total_sum <= total_sum + cache[3498];
endrule
rule s3500(sum_count == 3500);
  total_sum <= total_sum + cache[3499];
endrule
rule s3501(sum_count == 3501);
  total_sum <= total_sum + cache[3500];
endrule
rule s3502(sum_count == 3502);
  total_sum <= total_sum + cache[3501];
endrule
rule s3503(sum_count == 3503);
  total_sum <= total_sum + cache[3502];
endrule
rule s3504(sum_count == 3504);
  total_sum <= total_sum + cache[3503];
endrule
rule s3505(sum_count == 3505);
  total_sum <= total_sum + cache[3504];
endrule
rule s3506(sum_count == 3506);
  total_sum <= total_sum + cache[3505];
endrule
rule s3507(sum_count == 3507);
  total_sum <= total_sum + cache[3506];
endrule
rule s3508(sum_count == 3508);
  total_sum <= total_sum + cache[3507];
endrule
rule s3509(sum_count == 3509);
  total_sum <= total_sum + cache[3508];
endrule
rule s3510(sum_count == 3510);
  total_sum <= total_sum + cache[3509];
endrule
rule s3511(sum_count == 3511);
  total_sum <= total_sum + cache[3510];
endrule
rule s3512(sum_count == 3512);
  total_sum <= total_sum + cache[3511];
endrule
rule s3513(sum_count == 3513);
  total_sum <= total_sum + cache[3512];
endrule
rule s3514(sum_count == 3514);
  total_sum <= total_sum + cache[3513];
endrule
rule s3515(sum_count == 3515);
  total_sum <= total_sum + cache[3514];
endrule
rule s3516(sum_count == 3516);
  total_sum <= total_sum + cache[3515];
endrule
rule s3517(sum_count == 3517);
  total_sum <= total_sum + cache[3516];
endrule
rule s3518(sum_count == 3518);
  total_sum <= total_sum + cache[3517];
endrule
rule s3519(sum_count == 3519);
  total_sum <= total_sum + cache[3518];
endrule
rule s3520(sum_count == 3520);
  total_sum <= total_sum + cache[3519];
endrule
rule s3521(sum_count == 3521);
  total_sum <= total_sum + cache[3520];
endrule
rule s3522(sum_count == 3522);
  total_sum <= total_sum + cache[3521];
endrule
rule s3523(sum_count == 3523);
  total_sum <= total_sum + cache[3522];
endrule
rule s3524(sum_count == 3524);
  total_sum <= total_sum + cache[3523];
endrule
rule s3525(sum_count == 3525);
  total_sum <= total_sum + cache[3524];
endrule
rule s3526(sum_count == 3526);
  total_sum <= total_sum + cache[3525];
endrule
rule s3527(sum_count == 3527);
  total_sum <= total_sum + cache[3526];
endrule
rule s3528(sum_count == 3528);
  total_sum <= total_sum + cache[3527];
endrule
rule s3529(sum_count == 3529);
  total_sum <= total_sum + cache[3528];
endrule
rule s3530(sum_count == 3530);
  total_sum <= total_sum + cache[3529];
endrule
rule s3531(sum_count == 3531);
  total_sum <= total_sum + cache[3530];
endrule
rule s3532(sum_count == 3532);
  total_sum <= total_sum + cache[3531];
endrule
rule s3533(sum_count == 3533);
  total_sum <= total_sum + cache[3532];
endrule
rule s3534(sum_count == 3534);
  total_sum <= total_sum + cache[3533];
endrule
rule s3535(sum_count == 3535);
  total_sum <= total_sum + cache[3534];
endrule
rule s3536(sum_count == 3536);
  total_sum <= total_sum + cache[3535];
endrule
rule s3537(sum_count == 3537);
  total_sum <= total_sum + cache[3536];
endrule
rule s3538(sum_count == 3538);
  total_sum <= total_sum + cache[3537];
endrule
rule s3539(sum_count == 3539);
  total_sum <= total_sum + cache[3538];
endrule
rule s3540(sum_count == 3540);
  total_sum <= total_sum + cache[3539];
endrule
rule s3541(sum_count == 3541);
  total_sum <= total_sum + cache[3540];
endrule
rule s3542(sum_count == 3542);
  total_sum <= total_sum + cache[3541];
endrule
rule s3543(sum_count == 3543);
  total_sum <= total_sum + cache[3542];
endrule
rule s3544(sum_count == 3544);
  total_sum <= total_sum + cache[3543];
endrule
rule s3545(sum_count == 3545);
  total_sum <= total_sum + cache[3544];
endrule
rule s3546(sum_count == 3546);
  total_sum <= total_sum + cache[3545];
endrule
rule s3547(sum_count == 3547);
  total_sum <= total_sum + cache[3546];
endrule
rule s3548(sum_count == 3548);
  total_sum <= total_sum + cache[3547];
endrule
rule s3549(sum_count == 3549);
  total_sum <= total_sum + cache[3548];
endrule
rule s3550(sum_count == 3550);
  total_sum <= total_sum + cache[3549];
endrule
rule s3551(sum_count == 3551);
  total_sum <= total_sum + cache[3550];
endrule
rule s3552(sum_count == 3552);
  total_sum <= total_sum + cache[3551];
endrule
rule s3553(sum_count == 3553);
  total_sum <= total_sum + cache[3552];
endrule
rule s3554(sum_count == 3554);
  total_sum <= total_sum + cache[3553];
endrule
rule s3555(sum_count == 3555);
  total_sum <= total_sum + cache[3554];
endrule
rule s3556(sum_count == 3556);
  total_sum <= total_sum + cache[3555];
endrule
rule s3557(sum_count == 3557);
  total_sum <= total_sum + cache[3556];
endrule
rule s3558(sum_count == 3558);
  total_sum <= total_sum + cache[3557];
endrule
rule s3559(sum_count == 3559);
  total_sum <= total_sum + cache[3558];
endrule
rule s3560(sum_count == 3560);
  total_sum <= total_sum + cache[3559];
endrule
rule s3561(sum_count == 3561);
  total_sum <= total_sum + cache[3560];
endrule
rule s3562(sum_count == 3562);
  total_sum <= total_sum + cache[3561];
endrule
rule s3563(sum_count == 3563);
  total_sum <= total_sum + cache[3562];
endrule
rule s3564(sum_count == 3564);
  total_sum <= total_sum + cache[3563];
endrule
rule s3565(sum_count == 3565);
  total_sum <= total_sum + cache[3564];
endrule
rule s3566(sum_count == 3566);
  total_sum <= total_sum + cache[3565];
endrule
rule s3567(sum_count == 3567);
  total_sum <= total_sum + cache[3566];
endrule
rule s3568(sum_count == 3568);
  total_sum <= total_sum + cache[3567];
endrule
rule s3569(sum_count == 3569);
  total_sum <= total_sum + cache[3568];
endrule
rule s3570(sum_count == 3570);
  total_sum <= total_sum + cache[3569];
endrule
rule s3571(sum_count == 3571);
  total_sum <= total_sum + cache[3570];
endrule
rule s3572(sum_count == 3572);
  total_sum <= total_sum + cache[3571];
endrule
rule s3573(sum_count == 3573);
  total_sum <= total_sum + cache[3572];
endrule
rule s3574(sum_count == 3574);
  total_sum <= total_sum + cache[3573];
endrule
rule s3575(sum_count == 3575);
  total_sum <= total_sum + cache[3574];
endrule
rule s3576(sum_count == 3576);
  total_sum <= total_sum + cache[3575];
endrule
rule s3577(sum_count == 3577);
  total_sum <= total_sum + cache[3576];
endrule
rule s3578(sum_count == 3578);
  total_sum <= total_sum + cache[3577];
endrule
rule s3579(sum_count == 3579);
  total_sum <= total_sum + cache[3578];
endrule
rule s3580(sum_count == 3580);
  total_sum <= total_sum + cache[3579];
endrule
rule s3581(sum_count == 3581);
  total_sum <= total_sum + cache[3580];
endrule
rule s3582(sum_count == 3582);
  total_sum <= total_sum + cache[3581];
endrule
rule s3583(sum_count == 3583);
  total_sum <= total_sum + cache[3582];
endrule
rule s3584(sum_count == 3584);
  total_sum <= total_sum + cache[3583];
endrule
rule s3585(sum_count == 3585);
  total_sum <= total_sum + cache[3584];
endrule
rule s3586(sum_count == 3586);
  total_sum <= total_sum + cache[3585];
endrule
rule s3587(sum_count == 3587);
  total_sum <= total_sum + cache[3586];
endrule
rule s3588(sum_count == 3588);
  total_sum <= total_sum + cache[3587];
endrule
rule s3589(sum_count == 3589);
  total_sum <= total_sum + cache[3588];
endrule
rule s3590(sum_count == 3590);
  total_sum <= total_sum + cache[3589];
endrule
rule s3591(sum_count == 3591);
  total_sum <= total_sum + cache[3590];
endrule
rule s3592(sum_count == 3592);
  total_sum <= total_sum + cache[3591];
endrule
rule s3593(sum_count == 3593);
  total_sum <= total_sum + cache[3592];
endrule
rule s3594(sum_count == 3594);
  total_sum <= total_sum + cache[3593];
endrule
rule s3595(sum_count == 3595);
  total_sum <= total_sum + cache[3594];
endrule
rule s3596(sum_count == 3596);
  total_sum <= total_sum + cache[3595];
endrule
rule s3597(sum_count == 3597);
  total_sum <= total_sum + cache[3596];
endrule
rule s3598(sum_count == 3598);
  total_sum <= total_sum + cache[3597];
endrule
rule s3599(sum_count == 3599);
  total_sum <= total_sum + cache[3598];
endrule
rule s3600(sum_count == 3600);
  total_sum <= total_sum + cache[3599];
endrule
rule s3601(sum_count == 3601);
  total_sum <= total_sum + cache[3600];
endrule
rule s3602(sum_count == 3602);
  total_sum <= total_sum + cache[3601];
endrule
rule s3603(sum_count == 3603);
  total_sum <= total_sum + cache[3602];
endrule
rule s3604(sum_count == 3604);
  total_sum <= total_sum + cache[3603];
endrule
rule s3605(sum_count == 3605);
  total_sum <= total_sum + cache[3604];
endrule
rule s3606(sum_count == 3606);
  total_sum <= total_sum + cache[3605];
endrule
rule s3607(sum_count == 3607);
  total_sum <= total_sum + cache[3606];
endrule
rule s3608(sum_count == 3608);
  total_sum <= total_sum + cache[3607];
endrule
rule s3609(sum_count == 3609);
  total_sum <= total_sum + cache[3608];
endrule
rule s3610(sum_count == 3610);
  total_sum <= total_sum + cache[3609];
endrule
rule s3611(sum_count == 3611);
  total_sum <= total_sum + cache[3610];
endrule
rule s3612(sum_count == 3612);
  total_sum <= total_sum + cache[3611];
endrule
rule s3613(sum_count == 3613);
  total_sum <= total_sum + cache[3612];
endrule
rule s3614(sum_count == 3614);
  total_sum <= total_sum + cache[3613];
endrule
rule s3615(sum_count == 3615);
  total_sum <= total_sum + cache[3614];
endrule
rule s3616(sum_count == 3616);
  total_sum <= total_sum + cache[3615];
endrule
rule s3617(sum_count == 3617);
  total_sum <= total_sum + cache[3616];
endrule
rule s3618(sum_count == 3618);
  total_sum <= total_sum + cache[3617];
endrule
rule s3619(sum_count == 3619);
  total_sum <= total_sum + cache[3618];
endrule
rule s3620(sum_count == 3620);
  total_sum <= total_sum + cache[3619];
endrule
rule s3621(sum_count == 3621);
  total_sum <= total_sum + cache[3620];
endrule
rule s3622(sum_count == 3622);
  total_sum <= total_sum + cache[3621];
endrule
rule s3623(sum_count == 3623);
  total_sum <= total_sum + cache[3622];
endrule
rule s3624(sum_count == 3624);
  total_sum <= total_sum + cache[3623];
endrule
rule s3625(sum_count == 3625);
  total_sum <= total_sum + cache[3624];
endrule
rule s3626(sum_count == 3626);
  total_sum <= total_sum + cache[3625];
endrule
rule s3627(sum_count == 3627);
  total_sum <= total_sum + cache[3626];
endrule
rule s3628(sum_count == 3628);
  total_sum <= total_sum + cache[3627];
endrule
rule s3629(sum_count == 3629);
  total_sum <= total_sum + cache[3628];
endrule
rule s3630(sum_count == 3630);
  total_sum <= total_sum + cache[3629];
endrule
rule s3631(sum_count == 3631);
  total_sum <= total_sum + cache[3630];
endrule
rule s3632(sum_count == 3632);
  total_sum <= total_sum + cache[3631];
endrule
rule s3633(sum_count == 3633);
  total_sum <= total_sum + cache[3632];
endrule
rule s3634(sum_count == 3634);
  total_sum <= total_sum + cache[3633];
endrule
rule s3635(sum_count == 3635);
  total_sum <= total_sum + cache[3634];
endrule
rule s3636(sum_count == 3636);
  total_sum <= total_sum + cache[3635];
endrule
rule s3637(sum_count == 3637);
  total_sum <= total_sum + cache[3636];
endrule
rule s3638(sum_count == 3638);
  total_sum <= total_sum + cache[3637];
endrule
rule s3639(sum_count == 3639);
  total_sum <= total_sum + cache[3638];
endrule
rule s3640(sum_count == 3640);
  total_sum <= total_sum + cache[3639];
endrule
rule s3641(sum_count == 3641);
  total_sum <= total_sum + cache[3640];
endrule
rule s3642(sum_count == 3642);
  total_sum <= total_sum + cache[3641];
endrule
rule s3643(sum_count == 3643);
  total_sum <= total_sum + cache[3642];
endrule
rule s3644(sum_count == 3644);
  total_sum <= total_sum + cache[3643];
endrule
rule s3645(sum_count == 3645);
  total_sum <= total_sum + cache[3644];
endrule
rule s3646(sum_count == 3646);
  total_sum <= total_sum + cache[3645];
endrule
rule s3647(sum_count == 3647);
  total_sum <= total_sum + cache[3646];
endrule
rule s3648(sum_count == 3648);
  total_sum <= total_sum + cache[3647];
endrule
rule s3649(sum_count == 3649);
  total_sum <= total_sum + cache[3648];
endrule
rule s3650(sum_count == 3650);
  total_sum <= total_sum + cache[3649];
endrule
rule s3651(sum_count == 3651);
  total_sum <= total_sum + cache[3650];
endrule
rule s3652(sum_count == 3652);
  total_sum <= total_sum + cache[3651];
endrule
rule s3653(sum_count == 3653);
  total_sum <= total_sum + cache[3652];
endrule
rule s3654(sum_count == 3654);
  total_sum <= total_sum + cache[3653];
endrule
rule s3655(sum_count == 3655);
  total_sum <= total_sum + cache[3654];
endrule
rule s3656(sum_count == 3656);
  total_sum <= total_sum + cache[3655];
endrule
rule s3657(sum_count == 3657);
  total_sum <= total_sum + cache[3656];
endrule
rule s3658(sum_count == 3658);
  total_sum <= total_sum + cache[3657];
endrule
rule s3659(sum_count == 3659);
  total_sum <= total_sum + cache[3658];
endrule
rule s3660(sum_count == 3660);
  total_sum <= total_sum + cache[3659];
endrule
rule s3661(sum_count == 3661);
  total_sum <= total_sum + cache[3660];
endrule
rule s3662(sum_count == 3662);
  total_sum <= total_sum + cache[3661];
endrule
rule s3663(sum_count == 3663);
  total_sum <= total_sum + cache[3662];
endrule
rule s3664(sum_count == 3664);
  total_sum <= total_sum + cache[3663];
endrule
rule s3665(sum_count == 3665);
  total_sum <= total_sum + cache[3664];
endrule
rule s3666(sum_count == 3666);
  total_sum <= total_sum + cache[3665];
endrule
rule s3667(sum_count == 3667);
  total_sum <= total_sum + cache[3666];
endrule
rule s3668(sum_count == 3668);
  total_sum <= total_sum + cache[3667];
endrule
rule s3669(sum_count == 3669);
  total_sum <= total_sum + cache[3668];
endrule
rule s3670(sum_count == 3670);
  total_sum <= total_sum + cache[3669];
endrule
rule s3671(sum_count == 3671);
  total_sum <= total_sum + cache[3670];
endrule
rule s3672(sum_count == 3672);
  total_sum <= total_sum + cache[3671];
endrule
rule s3673(sum_count == 3673);
  total_sum <= total_sum + cache[3672];
endrule
rule s3674(sum_count == 3674);
  total_sum <= total_sum + cache[3673];
endrule
rule s3675(sum_count == 3675);
  total_sum <= total_sum + cache[3674];
endrule
rule s3676(sum_count == 3676);
  total_sum <= total_sum + cache[3675];
endrule
rule s3677(sum_count == 3677);
  total_sum <= total_sum + cache[3676];
endrule
rule s3678(sum_count == 3678);
  total_sum <= total_sum + cache[3677];
endrule
rule s3679(sum_count == 3679);
  total_sum <= total_sum + cache[3678];
endrule
rule s3680(sum_count == 3680);
  total_sum <= total_sum + cache[3679];
endrule
rule s3681(sum_count == 3681);
  total_sum <= total_sum + cache[3680];
endrule
rule s3682(sum_count == 3682);
  total_sum <= total_sum + cache[3681];
endrule
rule s3683(sum_count == 3683);
  total_sum <= total_sum + cache[3682];
endrule
rule s3684(sum_count == 3684);
  total_sum <= total_sum + cache[3683];
endrule
rule s3685(sum_count == 3685);
  total_sum <= total_sum + cache[3684];
endrule
rule s3686(sum_count == 3686);
  total_sum <= total_sum + cache[3685];
endrule
rule s3687(sum_count == 3687);
  total_sum <= total_sum + cache[3686];
endrule
rule s3688(sum_count == 3688);
  total_sum <= total_sum + cache[3687];
endrule
rule s3689(sum_count == 3689);
  total_sum <= total_sum + cache[3688];
endrule
rule s3690(sum_count == 3690);
  total_sum <= total_sum + cache[3689];
endrule
rule s3691(sum_count == 3691);
  total_sum <= total_sum + cache[3690];
endrule
rule s3692(sum_count == 3692);
  total_sum <= total_sum + cache[3691];
endrule
rule s3693(sum_count == 3693);
  total_sum <= total_sum + cache[3692];
endrule
rule s3694(sum_count == 3694);
  total_sum <= total_sum + cache[3693];
endrule
rule s3695(sum_count == 3695);
  total_sum <= total_sum + cache[3694];
endrule
rule s3696(sum_count == 3696);
  total_sum <= total_sum + cache[3695];
endrule
rule s3697(sum_count == 3697);
  total_sum <= total_sum + cache[3696];
endrule
rule s3698(sum_count == 3698);
  total_sum <= total_sum + cache[3697];
endrule
rule s3699(sum_count == 3699);
  total_sum <= total_sum + cache[3698];
endrule
rule s3700(sum_count == 3700);
  total_sum <= total_sum + cache[3699];
endrule
rule s3701(sum_count == 3701);
  total_sum <= total_sum + cache[3700];
endrule
rule s3702(sum_count == 3702);
  total_sum <= total_sum + cache[3701];
endrule
rule s3703(sum_count == 3703);
  total_sum <= total_sum + cache[3702];
endrule
rule s3704(sum_count == 3704);
  total_sum <= total_sum + cache[3703];
endrule
rule s3705(sum_count == 3705);
  total_sum <= total_sum + cache[3704];
endrule
rule s3706(sum_count == 3706);
  total_sum <= total_sum + cache[3705];
endrule
rule s3707(sum_count == 3707);
  total_sum <= total_sum + cache[3706];
endrule
rule s3708(sum_count == 3708);
  total_sum <= total_sum + cache[3707];
endrule
rule s3709(sum_count == 3709);
  total_sum <= total_sum + cache[3708];
endrule
rule s3710(sum_count == 3710);
  total_sum <= total_sum + cache[3709];
endrule
rule s3711(sum_count == 3711);
  total_sum <= total_sum + cache[3710];
endrule
rule s3712(sum_count == 3712);
  total_sum <= total_sum + cache[3711];
endrule
rule s3713(sum_count == 3713);
  total_sum <= total_sum + cache[3712];
endrule
rule s3714(sum_count == 3714);
  total_sum <= total_sum + cache[3713];
endrule
rule s3715(sum_count == 3715);
  total_sum <= total_sum + cache[3714];
endrule
rule s3716(sum_count == 3716);
  total_sum <= total_sum + cache[3715];
endrule
rule s3717(sum_count == 3717);
  total_sum <= total_sum + cache[3716];
endrule
rule s3718(sum_count == 3718);
  total_sum <= total_sum + cache[3717];
endrule
rule s3719(sum_count == 3719);
  total_sum <= total_sum + cache[3718];
endrule
rule s3720(sum_count == 3720);
  total_sum <= total_sum + cache[3719];
endrule
rule s3721(sum_count == 3721);
  total_sum <= total_sum + cache[3720];
endrule
rule s3722(sum_count == 3722);
  total_sum <= total_sum + cache[3721];
endrule
rule s3723(sum_count == 3723);
  total_sum <= total_sum + cache[3722];
endrule
rule s3724(sum_count == 3724);
  total_sum <= total_sum + cache[3723];
endrule
rule s3725(sum_count == 3725);
  total_sum <= total_sum + cache[3724];
endrule
rule s3726(sum_count == 3726);
  total_sum <= total_sum + cache[3725];
endrule
rule s3727(sum_count == 3727);
  total_sum <= total_sum + cache[3726];
endrule
rule s3728(sum_count == 3728);
  total_sum <= total_sum + cache[3727];
endrule
rule s3729(sum_count == 3729);
  total_sum <= total_sum + cache[3728];
endrule
rule s3730(sum_count == 3730);
  total_sum <= total_sum + cache[3729];
endrule
rule s3731(sum_count == 3731);
  total_sum <= total_sum + cache[3730];
endrule
rule s3732(sum_count == 3732);
  total_sum <= total_sum + cache[3731];
endrule
rule s3733(sum_count == 3733);
  total_sum <= total_sum + cache[3732];
endrule
rule s3734(sum_count == 3734);
  total_sum <= total_sum + cache[3733];
endrule
rule s3735(sum_count == 3735);
  total_sum <= total_sum + cache[3734];
endrule
rule s3736(sum_count == 3736);
  total_sum <= total_sum + cache[3735];
endrule
rule s3737(sum_count == 3737);
  total_sum <= total_sum + cache[3736];
endrule
rule s3738(sum_count == 3738);
  total_sum <= total_sum + cache[3737];
endrule
rule s3739(sum_count == 3739);
  total_sum <= total_sum + cache[3738];
endrule
rule s3740(sum_count == 3740);
  total_sum <= total_sum + cache[3739];
endrule
rule s3741(sum_count == 3741);
  total_sum <= total_sum + cache[3740];
endrule
rule s3742(sum_count == 3742);
  total_sum <= total_sum + cache[3741];
endrule
rule s3743(sum_count == 3743);
  total_sum <= total_sum + cache[3742];
endrule
rule s3744(sum_count == 3744);
  total_sum <= total_sum + cache[3743];
endrule
rule s3745(sum_count == 3745);
  total_sum <= total_sum + cache[3744];
endrule
rule s3746(sum_count == 3746);
  total_sum <= total_sum + cache[3745];
endrule
rule s3747(sum_count == 3747);
  total_sum <= total_sum + cache[3746];
endrule
rule s3748(sum_count == 3748);
  total_sum <= total_sum + cache[3747];
endrule
rule s3749(sum_count == 3749);
  total_sum <= total_sum + cache[3748];
endrule
rule s3750(sum_count == 3750);
  total_sum <= total_sum + cache[3749];
endrule
rule s3751(sum_count == 3751);
  total_sum <= total_sum + cache[3750];
endrule
rule s3752(sum_count == 3752);
  total_sum <= total_sum + cache[3751];
endrule
rule s3753(sum_count == 3753);
  total_sum <= total_sum + cache[3752];
endrule
rule s3754(sum_count == 3754);
  total_sum <= total_sum + cache[3753];
endrule
rule s3755(sum_count == 3755);
  total_sum <= total_sum + cache[3754];
endrule
rule s3756(sum_count == 3756);
  total_sum <= total_sum + cache[3755];
endrule
rule s3757(sum_count == 3757);
  total_sum <= total_sum + cache[3756];
endrule
rule s3758(sum_count == 3758);
  total_sum <= total_sum + cache[3757];
endrule
rule s3759(sum_count == 3759);
  total_sum <= total_sum + cache[3758];
endrule
rule s3760(sum_count == 3760);
  total_sum <= total_sum + cache[3759];
endrule
rule s3761(sum_count == 3761);
  total_sum <= total_sum + cache[3760];
endrule
rule s3762(sum_count == 3762);
  total_sum <= total_sum + cache[3761];
endrule
rule s3763(sum_count == 3763);
  total_sum <= total_sum + cache[3762];
endrule
rule s3764(sum_count == 3764);
  total_sum <= total_sum + cache[3763];
endrule
rule s3765(sum_count == 3765);
  total_sum <= total_sum + cache[3764];
endrule
rule s3766(sum_count == 3766);
  total_sum <= total_sum + cache[3765];
endrule
rule s3767(sum_count == 3767);
  total_sum <= total_sum + cache[3766];
endrule
rule s3768(sum_count == 3768);
  total_sum <= total_sum + cache[3767];
endrule
rule s3769(sum_count == 3769);
  total_sum <= total_sum + cache[3768];
endrule
rule s3770(sum_count == 3770);
  total_sum <= total_sum + cache[3769];
endrule
rule s3771(sum_count == 3771);
  total_sum <= total_sum + cache[3770];
endrule
rule s3772(sum_count == 3772);
  total_sum <= total_sum + cache[3771];
endrule
rule s3773(sum_count == 3773);
  total_sum <= total_sum + cache[3772];
endrule
rule s3774(sum_count == 3774);
  total_sum <= total_sum + cache[3773];
endrule
rule s3775(sum_count == 3775);
  total_sum <= total_sum + cache[3774];
endrule
rule s3776(sum_count == 3776);
  total_sum <= total_sum + cache[3775];
endrule
rule s3777(sum_count == 3777);
  total_sum <= total_sum + cache[3776];
endrule
rule s3778(sum_count == 3778);
  total_sum <= total_sum + cache[3777];
endrule
rule s3779(sum_count == 3779);
  total_sum <= total_sum + cache[3778];
endrule
rule s3780(sum_count == 3780);
  total_sum <= total_sum + cache[3779];
endrule
rule s3781(sum_count == 3781);
  total_sum <= total_sum + cache[3780];
endrule
rule s3782(sum_count == 3782);
  total_sum <= total_sum + cache[3781];
endrule
rule s3783(sum_count == 3783);
  total_sum <= total_sum + cache[3782];
endrule
rule s3784(sum_count == 3784);
  total_sum <= total_sum + cache[3783];
endrule
rule s3785(sum_count == 3785);
  total_sum <= total_sum + cache[3784];
endrule
rule s3786(sum_count == 3786);
  total_sum <= total_sum + cache[3785];
endrule
rule s3787(sum_count == 3787);
  total_sum <= total_sum + cache[3786];
endrule
rule s3788(sum_count == 3788);
  total_sum <= total_sum + cache[3787];
endrule
rule s3789(sum_count == 3789);
  total_sum <= total_sum + cache[3788];
endrule
rule s3790(sum_count == 3790);
  total_sum <= total_sum + cache[3789];
endrule
rule s3791(sum_count == 3791);
  total_sum <= total_sum + cache[3790];
endrule
rule s3792(sum_count == 3792);
  total_sum <= total_sum + cache[3791];
endrule
rule s3793(sum_count == 3793);
  total_sum <= total_sum + cache[3792];
endrule
rule s3794(sum_count == 3794);
  total_sum <= total_sum + cache[3793];
endrule
rule s3795(sum_count == 3795);
  total_sum <= total_sum + cache[3794];
endrule
rule s3796(sum_count == 3796);
  total_sum <= total_sum + cache[3795];
endrule
rule s3797(sum_count == 3797);
  total_sum <= total_sum + cache[3796];
endrule
rule s3798(sum_count == 3798);
  total_sum <= total_sum + cache[3797];
endrule
rule s3799(sum_count == 3799);
  total_sum <= total_sum + cache[3798];
endrule
rule s3800(sum_count == 3800);
  total_sum <= total_sum + cache[3799];
endrule
rule s3801(sum_count == 3801);
  total_sum <= total_sum + cache[3800];
endrule
rule s3802(sum_count == 3802);
  total_sum <= total_sum + cache[3801];
endrule
rule s3803(sum_count == 3803);
  total_sum <= total_sum + cache[3802];
endrule
rule s3804(sum_count == 3804);
  total_sum <= total_sum + cache[3803];
endrule
rule s3805(sum_count == 3805);
  total_sum <= total_sum + cache[3804];
endrule
rule s3806(sum_count == 3806);
  total_sum <= total_sum + cache[3805];
endrule
rule s3807(sum_count == 3807);
  total_sum <= total_sum + cache[3806];
endrule
rule s3808(sum_count == 3808);
  total_sum <= total_sum + cache[3807];
endrule
rule s3809(sum_count == 3809);
  total_sum <= total_sum + cache[3808];
endrule
rule s3810(sum_count == 3810);
  total_sum <= total_sum + cache[3809];
endrule
rule s3811(sum_count == 3811);
  total_sum <= total_sum + cache[3810];
endrule
rule s3812(sum_count == 3812);
  total_sum <= total_sum + cache[3811];
endrule
rule s3813(sum_count == 3813);
  total_sum <= total_sum + cache[3812];
endrule
rule s3814(sum_count == 3814);
  total_sum <= total_sum + cache[3813];
endrule
rule s3815(sum_count == 3815);
  total_sum <= total_sum + cache[3814];
endrule
rule s3816(sum_count == 3816);
  total_sum <= total_sum + cache[3815];
endrule
rule s3817(sum_count == 3817);
  total_sum <= total_sum + cache[3816];
endrule
rule s3818(sum_count == 3818);
  total_sum <= total_sum + cache[3817];
endrule
rule s3819(sum_count == 3819);
  total_sum <= total_sum + cache[3818];
endrule
rule s3820(sum_count == 3820);
  total_sum <= total_sum + cache[3819];
endrule
rule s3821(sum_count == 3821);
  total_sum <= total_sum + cache[3820];
endrule
rule s3822(sum_count == 3822);
  total_sum <= total_sum + cache[3821];
endrule
rule s3823(sum_count == 3823);
  total_sum <= total_sum + cache[3822];
endrule
rule s3824(sum_count == 3824);
  total_sum <= total_sum + cache[3823];
endrule
rule s3825(sum_count == 3825);
  total_sum <= total_sum + cache[3824];
endrule
rule s3826(sum_count == 3826);
  total_sum <= total_sum + cache[3825];
endrule
rule s3827(sum_count == 3827);
  total_sum <= total_sum + cache[3826];
endrule
rule s3828(sum_count == 3828);
  total_sum <= total_sum + cache[3827];
endrule
rule s3829(sum_count == 3829);
  total_sum <= total_sum + cache[3828];
endrule
rule s3830(sum_count == 3830);
  total_sum <= total_sum + cache[3829];
endrule
rule s3831(sum_count == 3831);
  total_sum <= total_sum + cache[3830];
endrule
rule s3832(sum_count == 3832);
  total_sum <= total_sum + cache[3831];
endrule
rule s3833(sum_count == 3833);
  total_sum <= total_sum + cache[3832];
endrule
rule s3834(sum_count == 3834);
  total_sum <= total_sum + cache[3833];
endrule
rule s3835(sum_count == 3835);
  total_sum <= total_sum + cache[3834];
endrule
rule s3836(sum_count == 3836);
  total_sum <= total_sum + cache[3835];
endrule
rule s3837(sum_count == 3837);
  total_sum <= total_sum + cache[3836];
endrule
rule s3838(sum_count == 3838);
  total_sum <= total_sum + cache[3837];
endrule
rule s3839(sum_count == 3839);
  total_sum <= total_sum + cache[3838];
endrule
rule s3840(sum_count == 3840);
  total_sum <= total_sum + cache[3839];
endrule
rule s3841(sum_count == 3841);
  total_sum <= total_sum + cache[3840];
endrule
rule s3842(sum_count == 3842);
  total_sum <= total_sum + cache[3841];
endrule
rule s3843(sum_count == 3843);
  total_sum <= total_sum + cache[3842];
endrule
rule s3844(sum_count == 3844);
  total_sum <= total_sum + cache[3843];
endrule
rule s3845(sum_count == 3845);
  total_sum <= total_sum + cache[3844];
endrule
rule s3846(sum_count == 3846);
  total_sum <= total_sum + cache[3845];
endrule
rule s3847(sum_count == 3847);
  total_sum <= total_sum + cache[3846];
endrule
rule s3848(sum_count == 3848);
  total_sum <= total_sum + cache[3847];
endrule
rule s3849(sum_count == 3849);
  total_sum <= total_sum + cache[3848];
endrule
rule s3850(sum_count == 3850);
  total_sum <= total_sum + cache[3849];
endrule
rule s3851(sum_count == 3851);
  total_sum <= total_sum + cache[3850];
endrule
rule s3852(sum_count == 3852);
  total_sum <= total_sum + cache[3851];
endrule
rule s3853(sum_count == 3853);
  total_sum <= total_sum + cache[3852];
endrule
rule s3854(sum_count == 3854);
  total_sum <= total_sum + cache[3853];
endrule
rule s3855(sum_count == 3855);
  total_sum <= total_sum + cache[3854];
endrule
rule s3856(sum_count == 3856);
  total_sum <= total_sum + cache[3855];
endrule
rule s3857(sum_count == 3857);
  total_sum <= total_sum + cache[3856];
endrule
rule s3858(sum_count == 3858);
  total_sum <= total_sum + cache[3857];
endrule
rule s3859(sum_count == 3859);
  total_sum <= total_sum + cache[3858];
endrule
rule s3860(sum_count == 3860);
  total_sum <= total_sum + cache[3859];
endrule
rule s3861(sum_count == 3861);
  total_sum <= total_sum + cache[3860];
endrule
rule s3862(sum_count == 3862);
  total_sum <= total_sum + cache[3861];
endrule
rule s3863(sum_count == 3863);
  total_sum <= total_sum + cache[3862];
endrule
rule s3864(sum_count == 3864);
  total_sum <= total_sum + cache[3863];
endrule
rule s3865(sum_count == 3865);
  total_sum <= total_sum + cache[3864];
endrule
rule s3866(sum_count == 3866);
  total_sum <= total_sum + cache[3865];
endrule
rule s3867(sum_count == 3867);
  total_sum <= total_sum + cache[3866];
endrule
rule s3868(sum_count == 3868);
  total_sum <= total_sum + cache[3867];
endrule
rule s3869(sum_count == 3869);
  total_sum <= total_sum + cache[3868];
endrule
rule s3870(sum_count == 3870);
  total_sum <= total_sum + cache[3869];
endrule
rule s3871(sum_count == 3871);
  total_sum <= total_sum + cache[3870];
endrule
rule s3872(sum_count == 3872);
  total_sum <= total_sum + cache[3871];
endrule
rule s3873(sum_count == 3873);
  total_sum <= total_sum + cache[3872];
endrule
rule s3874(sum_count == 3874);
  total_sum <= total_sum + cache[3873];
endrule
rule s3875(sum_count == 3875);
  total_sum <= total_sum + cache[3874];
endrule
rule s3876(sum_count == 3876);
  total_sum <= total_sum + cache[3875];
endrule
rule s3877(sum_count == 3877);
  total_sum <= total_sum + cache[3876];
endrule
rule s3878(sum_count == 3878);
  total_sum <= total_sum + cache[3877];
endrule
rule s3879(sum_count == 3879);
  total_sum <= total_sum + cache[3878];
endrule
rule s3880(sum_count == 3880);
  total_sum <= total_sum + cache[3879];
endrule
rule s3881(sum_count == 3881);
  total_sum <= total_sum + cache[3880];
endrule
rule s3882(sum_count == 3882);
  total_sum <= total_sum + cache[3881];
endrule
rule s3883(sum_count == 3883);
  total_sum <= total_sum + cache[3882];
endrule
rule s3884(sum_count == 3884);
  total_sum <= total_sum + cache[3883];
endrule
rule s3885(sum_count == 3885);
  total_sum <= total_sum + cache[3884];
endrule
rule s3886(sum_count == 3886);
  total_sum <= total_sum + cache[3885];
endrule
rule s3887(sum_count == 3887);
  total_sum <= total_sum + cache[3886];
endrule
rule s3888(sum_count == 3888);
  total_sum <= total_sum + cache[3887];
endrule
rule s3889(sum_count == 3889);
  total_sum <= total_sum + cache[3888];
endrule
rule s3890(sum_count == 3890);
  total_sum <= total_sum + cache[3889];
endrule
rule s3891(sum_count == 3891);
  total_sum <= total_sum + cache[3890];
endrule
rule s3892(sum_count == 3892);
  total_sum <= total_sum + cache[3891];
endrule
rule s3893(sum_count == 3893);
  total_sum <= total_sum + cache[3892];
endrule
rule s3894(sum_count == 3894);
  total_sum <= total_sum + cache[3893];
endrule
rule s3895(sum_count == 3895);
  total_sum <= total_sum + cache[3894];
endrule
rule s3896(sum_count == 3896);
  total_sum <= total_sum + cache[3895];
endrule
rule s3897(sum_count == 3897);
  total_sum <= total_sum + cache[3896];
endrule
rule s3898(sum_count == 3898);
  total_sum <= total_sum + cache[3897];
endrule
rule s3899(sum_count == 3899);
  total_sum <= total_sum + cache[3898];
endrule
rule s3900(sum_count == 3900);
  total_sum <= total_sum + cache[3899];
endrule
rule s3901(sum_count == 3901);
  total_sum <= total_sum + cache[3900];
endrule
rule s3902(sum_count == 3902);
  total_sum <= total_sum + cache[3901];
endrule
rule s3903(sum_count == 3903);
  total_sum <= total_sum + cache[3902];
endrule
rule s3904(sum_count == 3904);
  total_sum <= total_sum + cache[3903];
endrule
rule s3905(sum_count == 3905);
  total_sum <= total_sum + cache[3904];
endrule
rule s3906(sum_count == 3906);
  total_sum <= total_sum + cache[3905];
endrule
rule s3907(sum_count == 3907);
  total_sum <= total_sum + cache[3906];
endrule
rule s3908(sum_count == 3908);
  total_sum <= total_sum + cache[3907];
endrule
rule s3909(sum_count == 3909);
  total_sum <= total_sum + cache[3908];
endrule
rule s3910(sum_count == 3910);
  total_sum <= total_sum + cache[3909];
endrule
rule s3911(sum_count == 3911);
  total_sum <= total_sum + cache[3910];
endrule
rule s3912(sum_count == 3912);
  total_sum <= total_sum + cache[3911];
endrule
rule s3913(sum_count == 3913);
  total_sum <= total_sum + cache[3912];
endrule
rule s3914(sum_count == 3914);
  total_sum <= total_sum + cache[3913];
endrule
rule s3915(sum_count == 3915);
  total_sum <= total_sum + cache[3914];
endrule
rule s3916(sum_count == 3916);
  total_sum <= total_sum + cache[3915];
endrule
rule s3917(sum_count == 3917);
  total_sum <= total_sum + cache[3916];
endrule
rule s3918(sum_count == 3918);
  total_sum <= total_sum + cache[3917];
endrule
rule s3919(sum_count == 3919);
  total_sum <= total_sum + cache[3918];
endrule
rule s3920(sum_count == 3920);
  total_sum <= total_sum + cache[3919];
endrule
rule s3921(sum_count == 3921);
  total_sum <= total_sum + cache[3920];
endrule
rule s3922(sum_count == 3922);
  total_sum <= total_sum + cache[3921];
endrule
rule s3923(sum_count == 3923);
  total_sum <= total_sum + cache[3922];
endrule
rule s3924(sum_count == 3924);
  total_sum <= total_sum + cache[3923];
endrule
rule s3925(sum_count == 3925);
  total_sum <= total_sum + cache[3924];
endrule
rule s3926(sum_count == 3926);
  total_sum <= total_sum + cache[3925];
endrule
rule s3927(sum_count == 3927);
  total_sum <= total_sum + cache[3926];
endrule
rule s3928(sum_count == 3928);
  total_sum <= total_sum + cache[3927];
endrule
rule s3929(sum_count == 3929);
  total_sum <= total_sum + cache[3928];
endrule
rule s3930(sum_count == 3930);
  total_sum <= total_sum + cache[3929];
endrule
rule s3931(sum_count == 3931);
  total_sum <= total_sum + cache[3930];
endrule
rule s3932(sum_count == 3932);
  total_sum <= total_sum + cache[3931];
endrule
rule s3933(sum_count == 3933);
  total_sum <= total_sum + cache[3932];
endrule
rule s3934(sum_count == 3934);
  total_sum <= total_sum + cache[3933];
endrule
rule s3935(sum_count == 3935);
  total_sum <= total_sum + cache[3934];
endrule
rule s3936(sum_count == 3936);
  total_sum <= total_sum + cache[3935];
endrule
rule s3937(sum_count == 3937);
  total_sum <= total_sum + cache[3936];
endrule
rule s3938(sum_count == 3938);
  total_sum <= total_sum + cache[3937];
endrule
rule s3939(sum_count == 3939);
  total_sum <= total_sum + cache[3938];
endrule
rule s3940(sum_count == 3940);
  total_sum <= total_sum + cache[3939];
endrule
rule s3941(sum_count == 3941);
  total_sum <= total_sum + cache[3940];
endrule
rule s3942(sum_count == 3942);
  total_sum <= total_sum + cache[3941];
endrule
rule s3943(sum_count == 3943);
  total_sum <= total_sum + cache[3942];
endrule
rule s3944(sum_count == 3944);
  total_sum <= total_sum + cache[3943];
endrule
rule s3945(sum_count == 3945);
  total_sum <= total_sum + cache[3944];
endrule
rule s3946(sum_count == 3946);
  total_sum <= total_sum + cache[3945];
endrule
rule s3947(sum_count == 3947);
  total_sum <= total_sum + cache[3946];
endrule
rule s3948(sum_count == 3948);
  total_sum <= total_sum + cache[3947];
endrule
rule s3949(sum_count == 3949);
  total_sum <= total_sum + cache[3948];
endrule
rule s3950(sum_count == 3950);
  total_sum <= total_sum + cache[3949];
endrule
rule s3951(sum_count == 3951);
  total_sum <= total_sum + cache[3950];
endrule
rule s3952(sum_count == 3952);
  total_sum <= total_sum + cache[3951];
endrule
rule s3953(sum_count == 3953);
  total_sum <= total_sum + cache[3952];
endrule
rule s3954(sum_count == 3954);
  total_sum <= total_sum + cache[3953];
endrule
rule s3955(sum_count == 3955);
  total_sum <= total_sum + cache[3954];
endrule
rule s3956(sum_count == 3956);
  total_sum <= total_sum + cache[3955];
endrule
rule s3957(sum_count == 3957);
  total_sum <= total_sum + cache[3956];
endrule
rule s3958(sum_count == 3958);
  total_sum <= total_sum + cache[3957];
endrule
rule s3959(sum_count == 3959);
  total_sum <= total_sum + cache[3958];
endrule
rule s3960(sum_count == 3960);
  total_sum <= total_sum + cache[3959];
endrule
rule s3961(sum_count == 3961);
  total_sum <= total_sum + cache[3960];
endrule
rule s3962(sum_count == 3962);
  total_sum <= total_sum + cache[3961];
endrule
rule s3963(sum_count == 3963);
  total_sum <= total_sum + cache[3962];
endrule
rule s3964(sum_count == 3964);
  total_sum <= total_sum + cache[3963];
endrule
rule s3965(sum_count == 3965);
  total_sum <= total_sum + cache[3964];
endrule
rule s3966(sum_count == 3966);
  total_sum <= total_sum + cache[3965];
endrule
rule s3967(sum_count == 3967);
  total_sum <= total_sum + cache[3966];
endrule
rule s3968(sum_count == 3968);
  total_sum <= total_sum + cache[3967];
endrule
rule s3969(sum_count == 3969);
  total_sum <= total_sum + cache[3968];
endrule
rule s3970(sum_count == 3970);
  total_sum <= total_sum + cache[3969];
endrule
rule s3971(sum_count == 3971);
  total_sum <= total_sum + cache[3970];
endrule
rule s3972(sum_count == 3972);
  total_sum <= total_sum + cache[3971];
endrule
rule s3973(sum_count == 3973);
  total_sum <= total_sum + cache[3972];
endrule
rule s3974(sum_count == 3974);
  total_sum <= total_sum + cache[3973];
endrule
rule s3975(sum_count == 3975);
  total_sum <= total_sum + cache[3974];
endrule
rule s3976(sum_count == 3976);
  total_sum <= total_sum + cache[3975];
endrule
rule s3977(sum_count == 3977);
  total_sum <= total_sum + cache[3976];
endrule
rule s3978(sum_count == 3978);
  total_sum <= total_sum + cache[3977];
endrule
rule s3979(sum_count == 3979);
  total_sum <= total_sum + cache[3978];
endrule
rule s3980(sum_count == 3980);
  total_sum <= total_sum + cache[3979];
endrule
rule s3981(sum_count == 3981);
  total_sum <= total_sum + cache[3980];
endrule
rule s3982(sum_count == 3982);
  total_sum <= total_sum + cache[3981];
endrule
rule s3983(sum_count == 3983);
  total_sum <= total_sum + cache[3982];
endrule
rule s3984(sum_count == 3984);
  total_sum <= total_sum + cache[3983];
endrule
rule s3985(sum_count == 3985);
  total_sum <= total_sum + cache[3984];
endrule
rule s3986(sum_count == 3986);
  total_sum <= total_sum + cache[3985];
endrule
rule s3987(sum_count == 3987);
  total_sum <= total_sum + cache[3986];
endrule
rule s3988(sum_count == 3988);
  total_sum <= total_sum + cache[3987];
endrule
rule s3989(sum_count == 3989);
  total_sum <= total_sum + cache[3988];
endrule
rule s3990(sum_count == 3990);
  total_sum <= total_sum + cache[3989];
endrule
rule s3991(sum_count == 3991);
  total_sum <= total_sum + cache[3990];
endrule
rule s3992(sum_count == 3992);
  total_sum <= total_sum + cache[3991];
endrule
rule s3993(sum_count == 3993);
  total_sum <= total_sum + cache[3992];
endrule
rule s3994(sum_count == 3994);
  total_sum <= total_sum + cache[3993];
endrule
rule s3995(sum_count == 3995);
  total_sum <= total_sum + cache[3994];
endrule
rule s3996(sum_count == 3996);
  total_sum <= total_sum + cache[3995];
endrule
rule s3997(sum_count == 3997);
  total_sum <= total_sum + cache[3996];
endrule
rule s3998(sum_count == 3998);
  total_sum <= total_sum + cache[3997];
endrule
rule s3999(sum_count == 3999);
  total_sum <= total_sum + cache[3998];
endrule
rule s4000(sum_count == 4000);
  total_sum <= total_sum + cache[3999];
endrule
rule s4001(sum_count == 4001);
  total_sum <= total_sum + cache[4000];
endrule
rule s4002(sum_count == 4002);
  total_sum <= total_sum + cache[4001];
endrule
rule s4003(sum_count == 4003);
  total_sum <= total_sum + cache[4002];
endrule
rule s4004(sum_count == 4004);
  total_sum <= total_sum + cache[4003];
endrule
rule s4005(sum_count == 4005);
  total_sum <= total_sum + cache[4004];
endrule
rule s4006(sum_count == 4006);
  total_sum <= total_sum + cache[4005];
endrule
rule s4007(sum_count == 4007);
  total_sum <= total_sum + cache[4006];
endrule
rule s4008(sum_count == 4008);
  total_sum <= total_sum + cache[4007];
endrule
rule s4009(sum_count == 4009);
  total_sum <= total_sum + cache[4008];
endrule
rule s4010(sum_count == 4010);
  total_sum <= total_sum + cache[4009];
endrule
rule s4011(sum_count == 4011);
  total_sum <= total_sum + cache[4010];
endrule
rule s4012(sum_count == 4012);
  total_sum <= total_sum + cache[4011];
endrule
rule s4013(sum_count == 4013);
  total_sum <= total_sum + cache[4012];
endrule
rule s4014(sum_count == 4014);
  total_sum <= total_sum + cache[4013];
endrule
rule s4015(sum_count == 4015);
  total_sum <= total_sum + cache[4014];
endrule
rule s4016(sum_count == 4016);
  total_sum <= total_sum + cache[4015];
endrule
rule s4017(sum_count == 4017);
  total_sum <= total_sum + cache[4016];
endrule
rule s4018(sum_count == 4018);
  total_sum <= total_sum + cache[4017];
endrule
rule s4019(sum_count == 4019);
  total_sum <= total_sum + cache[4018];
endrule
rule s4020(sum_count == 4020);
  total_sum <= total_sum + cache[4019];
endrule
rule s4021(sum_count == 4021);
  total_sum <= total_sum + cache[4020];
endrule
rule s4022(sum_count == 4022);
  total_sum <= total_sum + cache[4021];
endrule
rule s4023(sum_count == 4023);
  total_sum <= total_sum + cache[4022];
endrule
rule s4024(sum_count == 4024);
  total_sum <= total_sum + cache[4023];
endrule
rule s4025(sum_count == 4025);
  total_sum <= total_sum + cache[4024];
endrule
rule s4026(sum_count == 4026);
  total_sum <= total_sum + cache[4025];
endrule
rule s4027(sum_count == 4027);
  total_sum <= total_sum + cache[4026];
endrule
rule s4028(sum_count == 4028);
  total_sum <= total_sum + cache[4027];
endrule
rule s4029(sum_count == 4029);
  total_sum <= total_sum + cache[4028];
endrule
rule s4030(sum_count == 4030);
  total_sum <= total_sum + cache[4029];
endrule
rule s4031(sum_count == 4031);
  total_sum <= total_sum + cache[4030];
endrule
rule s4032(sum_count == 4032);
  total_sum <= total_sum + cache[4031];
endrule
rule s4033(sum_count == 4033);
  total_sum <= total_sum + cache[4032];
endrule
rule s4034(sum_count == 4034);
  total_sum <= total_sum + cache[4033];
endrule
rule s4035(sum_count == 4035);
  total_sum <= total_sum + cache[4034];
endrule
rule s4036(sum_count == 4036);
  total_sum <= total_sum + cache[4035];
endrule
rule s4037(sum_count == 4037);
  total_sum <= total_sum + cache[4036];
endrule
rule s4038(sum_count == 4038);
  total_sum <= total_sum + cache[4037];
endrule
rule s4039(sum_count == 4039);
  total_sum <= total_sum + cache[4038];
endrule
rule s4040(sum_count == 4040);
  total_sum <= total_sum + cache[4039];
endrule
rule s4041(sum_count == 4041);
  total_sum <= total_sum + cache[4040];
endrule
rule s4042(sum_count == 4042);
  total_sum <= total_sum + cache[4041];
endrule
rule s4043(sum_count == 4043);
  total_sum <= total_sum + cache[4042];
endrule
rule s4044(sum_count == 4044);
  total_sum <= total_sum + cache[4043];
endrule
rule s4045(sum_count == 4045);
  total_sum <= total_sum + cache[4044];
endrule
rule s4046(sum_count == 4046);
  total_sum <= total_sum + cache[4045];
endrule
rule s4047(sum_count == 4047);
  total_sum <= total_sum + cache[4046];
endrule
rule s4048(sum_count == 4048);
  total_sum <= total_sum + cache[4047];
endrule
rule s4049(sum_count == 4049);
  total_sum <= total_sum + cache[4048];
endrule
rule s4050(sum_count == 4050);
  total_sum <= total_sum + cache[4049];
endrule
rule s4051(sum_count == 4051);
  total_sum <= total_sum + cache[4050];
endrule
rule s4052(sum_count == 4052);
  total_sum <= total_sum + cache[4051];
endrule
rule s4053(sum_count == 4053);
  total_sum <= total_sum + cache[4052];
endrule
rule s4054(sum_count == 4054);
  total_sum <= total_sum + cache[4053];
endrule
rule s4055(sum_count == 4055);
  total_sum <= total_sum + cache[4054];
endrule
rule s4056(sum_count == 4056);
  total_sum <= total_sum + cache[4055];
endrule
rule s4057(sum_count == 4057);
  total_sum <= total_sum + cache[4056];
endrule
rule s4058(sum_count == 4058);
  total_sum <= total_sum + cache[4057];
endrule
rule s4059(sum_count == 4059);
  total_sum <= total_sum + cache[4058];
endrule
rule s4060(sum_count == 4060);
  total_sum <= total_sum + cache[4059];
endrule
rule s4061(sum_count == 4061);
  total_sum <= total_sum + cache[4060];
endrule
rule s4062(sum_count == 4062);
  total_sum <= total_sum + cache[4061];
endrule
rule s4063(sum_count == 4063);
  total_sum <= total_sum + cache[4062];
endrule
rule s4064(sum_count == 4064);
  total_sum <= total_sum + cache[4063];
endrule
rule s4065(sum_count == 4065);
  total_sum <= total_sum + cache[4064];
endrule
rule s4066(sum_count == 4066);
  total_sum <= total_sum + cache[4065];
endrule
rule s4067(sum_count == 4067);
  total_sum <= total_sum + cache[4066];
endrule
rule s4068(sum_count == 4068);
  total_sum <= total_sum + cache[4067];
endrule
rule s4069(sum_count == 4069);
  total_sum <= total_sum + cache[4068];
endrule
rule s4070(sum_count == 4070);
  total_sum <= total_sum + cache[4069];
endrule
rule s4071(sum_count == 4071);
  total_sum <= total_sum + cache[4070];
endrule
rule s4072(sum_count == 4072);
  total_sum <= total_sum + cache[4071];
endrule
rule s4073(sum_count == 4073);
  total_sum <= total_sum + cache[4072];
endrule
rule s4074(sum_count == 4074);
  total_sum <= total_sum + cache[4073];
endrule
rule s4075(sum_count == 4075);
  total_sum <= total_sum + cache[4074];
endrule
rule s4076(sum_count == 4076);
  total_sum <= total_sum + cache[4075];
endrule
rule s4077(sum_count == 4077);
  total_sum <= total_sum + cache[4076];
endrule
rule s4078(sum_count == 4078);
  total_sum <= total_sum + cache[4077];
endrule
rule s4079(sum_count == 4079);
  total_sum <= total_sum + cache[4078];
endrule
rule s4080(sum_count == 4080);
  total_sum <= total_sum + cache[4079];
endrule
rule s4081(sum_count == 4081);
  total_sum <= total_sum + cache[4080];
endrule
rule s4082(sum_count == 4082);
  total_sum <= total_sum + cache[4081];
endrule
rule s4083(sum_count == 4083);
  total_sum <= total_sum + cache[4082];
endrule
rule s4084(sum_count == 4084);
  total_sum <= total_sum + cache[4083];
endrule
rule s4085(sum_count == 4085);
  total_sum <= total_sum + cache[4084];
endrule
rule s4086(sum_count == 4086);
  total_sum <= total_sum + cache[4085];
endrule
rule s4087(sum_count == 4087);
  total_sum <= total_sum + cache[4086];
endrule
rule s4088(sum_count == 4088);
  total_sum <= total_sum + cache[4087];
endrule
rule s4089(sum_count == 4089);
  total_sum <= total_sum + cache[4088];
endrule
rule s4090(sum_count == 4090);
  total_sum <= total_sum + cache[4089];
endrule
rule s4091(sum_count == 4091);
  total_sum <= total_sum + cache[4090];
endrule
rule s4092(sum_count == 4092);
  total_sum <= total_sum + cache[4091];
endrule
rule s4093(sum_count == 4093);
  total_sum <= total_sum + cache[4092];
endrule
rule s4094(sum_count == 4094);
  total_sum <= total_sum + cache[4093];
endrule
rule s4095(sum_count == 4095);
  total_sum <= total_sum + cache[4094];
endrule
rule s4096(sum_count == 4096);
  total_sum <= total_sum + cache[4095];
endrule
        method Action put(DataType datas) if(ent < L0);
                      Bit#(MEMWORD) x = zeroExtend(pack(datas));
                      inQ <= (inQ << 8) | x;
                      ent <= ent + 1;
                  endmethod


        method Bit#(16) get;
                return pack(total_sum);
        endmethod
endmodule
endpackage